
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY voltage2distance IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      distance       :  OUT   STD_LOGIC_VECTOR(12 DOWNTO 0));  
END voltage2distance;

ARCHITECTURE behavior OF voltage2distance IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	4095	)	,
(	3299	)	,
(	3299	)	,
(	3299	)	,
(	3299	)	,
(	3294	)	,
(	3288	)	,
(	3282	)	,
(	3276	)	,
(	3270	)	,
(	3264	)	,
(	3258	)	,
(	3252	)	,
(	3246	)	,
(	3240	)	,
(	3234	)	,
(	3228	)	,
(	3222	)	,
(	3216	)	,
(	3210	)	,
(	3204	)	,
(	3198	)	,
(	3192	)	,
(	3186	)	,
(	3180	)	,
(	3174	)	,
(	3168	)	,
(	3162	)	,
(	3157	)	,
(	3151	)	,
(	3145	)	,
(	3139	)	,
(	3133	)	,
(	3127	)	,
(	3122	)	,
(	3116	)	,
(	3110	)	,
(	3104	)	,
(	3099	)	,
(	3093	)	,
(	3087	)	,
(	3082	)	,
(	3076	)	,
(	3070	)	,
(	3064	)	,
(	3059	)	,
(	3053	)	,
(	3048	)	,
(	3042	)	,
(	3036	)	,
(	3031	)	,
(	3025	)	,
(	3020	)	,
(	3014	)	,
(	3008	)	,
(	3003	)	,
(	2997	)	,
(	2992	)	,
(	2986	)	,
(	2981	)	,
(	2975	)	,
(	2970	)	,
(	2964	)	,
(	2959	)	,
(	2953	)	,
(	2948	)	,
(	2943	)	,
(	2937	)	,
(	2932	)	,
(	2926	)	,
(	2921	)	,
(	2916	)	,
(	2910	)	,
(	2905	)	,
(	2900	)	,
(	2894	)	,
(	2889	)	,
(	2884	)	,
(	2878	)	,
(	2873	)	,
(	2868	)	,
(	2863	)	,
(	2857	)	,
(	2852	)	,
(	2847	)	,
(	2842	)	,
(	2836	)	,
(	2831	)	,
(	2826	)	,
(	2821	)	,
(	2816	)	,
(	2811	)	,
(	2805	)	,
(	2800	)	,
(	2795	)	,
(	2790	)	,
(	2785	)	,
(	2780	)	,
(	2775	)	,
(	2770	)	,
(	2765	)	,
(	2760	)	,
(	2755	)	,
(	2750	)	,
(	2745	)	,
(	2740	)	,
(	2735	)	,
(	2730	)	,
(	2725	)	,
(	2720	)	,
(	2715	)	,
(	2710	)	,
(	2705	)	,
(	2700	)	,
(	2695	)	,
(	2690	)	,
(	2685	)	,
(	2680	)	,
(	2675	)	,
(	2671	)	,
(	2666	)	,
(	2661	)	,
(	2656	)	,
(	2651	)	,
(	2646	)	,
(	2642	)	,
(	2637	)	,
(	2632	)	,
(	2627	)	,
(	2622	)	,
(	2618	)	,
(	2613	)	,
(	2608	)	,
(	2603	)	,
(	2599	)	,
(	2594	)	,
(	2589	)	,
(	2585	)	,
(	2580	)	,
(	2575	)	,
(	2571	)	,
(	2566	)	,
(	2561	)	,
(	2557	)	,
(	2552	)	,
(	2548	)	,
(	2543	)	,
(	2538	)	,
(	2534	)	,
(	2529	)	,
(	2525	)	,
(	2520	)	,
(	2516	)	,
(	2511	)	,
(	2507	)	,
(	2502	)	,
(	2498	)	,
(	2493	)	,
(	2489	)	,
(	2484	)	,
(	2480	)	,
(	2475	)	,
(	2471	)	,
(	2466	)	,
(	2462	)	,
(	2458	)	,
(	2453	)	,
(	2449	)	,
(	2444	)	,
(	2440	)	,
(	2436	)	,
(	2431	)	,
(	2427	)	,
(	2423	)	,
(	2418	)	,
(	2414	)	,
(	2410	)	,
(	2405	)	,
(	2401	)	,
(	2397	)	,
(	2392	)	,
(	2388	)	,
(	2384	)	,
(	2380	)	,
(	2375	)	,
(	2371	)	,
(	2367	)	,
(	2363	)	,
(	2359	)	,
(	2354	)	,
(	2350	)	,
(	2346	)	,
(	2342	)	,
(	2338	)	,
(	2334	)	,
(	2330	)	,
(	2325	)	,
(	2321	)	,
(	2317	)	,
(	2313	)	,
(	2309	)	,
(	2305	)	,
(	2301	)	,
(	2297	)	,
(	2293	)	,
(	2289	)	,
(	2285	)	,
(	2281	)	,
(	2277	)	,
(	2273	)	,
(	2269	)	,
(	2265	)	,
(	2261	)	,
(	2257	)	,
(	2253	)	,
(	2249	)	,
(	2245	)	,
(	2241	)	,
(	2237	)	,
(	2233	)	,
(	2229	)	,
(	2225	)	,
(	2221	)	,
(	2217	)	,
(	2214	)	,
(	2210	)	,
(	2206	)	,
(	2202	)	,
(	2198	)	,
(	2194	)	,
(	2190	)	,
(	2187	)	,
(	2183	)	,
(	2179	)	,
(	2175	)	,
(	2171	)	,
(	2168	)	,
(	2164	)	,
(	2160	)	,
(	2156	)	,
(	2153	)	,
(	2149	)	,
(	2145	)	,
(	2141	)	,
(	2138	)	,
(	2134	)	,
(	2130	)	,
(	2127	)	,
(	2123	)	,
(	2119	)	,
(	2116	)	,
(	2112	)	,
(	2108	)	,
(	2105	)	,
(	2101	)	,
(	2098	)	,
(	2094	)	,
(	2090	)	,
(	2087	)	,
(	2083	)	,
(	2080	)	,
(	2076	)	,
(	2072	)	,
(	2069	)	,
(	2065	)	,
(	2062	)	,
(	2058	)	,
(	2055	)	,
(	2051	)	,
(	2048	)	,
(	2044	)	,
(	2041	)	,
(	2037	)	,
(	2034	)	,
(	2030	)	,
(	2027	)	,
(	2023	)	,
(	2020	)	,
(	2017	)	,
(	2013	)	,
(	2010	)	,
(	2006	)	,
(	2003	)	,
(	2000	)	,
(	1996	)	,
(	1993	)	,
(	1989	)	,
(	1986	)	,
(	1983	)	,
(	1979	)	,
(	1976	)	,
(	1973	)	,
(	1969	)	,
(	1966	)	,
(	1963	)	,
(	1959	)	,
(	1956	)	,
(	1953	)	,
(	1950	)	,
(	1946	)	,
(	1943	)	,
(	1940	)	,
(	1937	)	,
(	1933	)	,
(	1930	)	,
(	1927	)	,
(	1924	)	,
(	1920	)	,
(	1917	)	,
(	1914	)	,
(	1911	)	,
(	1908	)	,
(	1905	)	,
(	1901	)	,
(	1898	)	,
(	1895	)	,
(	1892	)	,
(	1889	)	,
(	1886	)	,
(	1883	)	,
(	1879	)	,
(	1876	)	,
(	1873	)	,
(	1870	)	,
(	1867	)	,
(	1864	)	,
(	1861	)	,
(	1858	)	,
(	1855	)	,
(	1852	)	,
(	1849	)	,
(	1846	)	,
(	1843	)	,
(	1840	)	,
(	1837	)	,
(	1834	)	,
(	1831	)	,
(	1828	)	,
(	1825	)	,
(	1822	)	,
(	1819	)	,
(	1816	)	,
(	1813	)	,
(	1810	)	,
(	1807	)	,
(	1804	)	,
(	1801	)	,
(	1798	)	,
(	1795	)	,
(	1792	)	,
(	1790	)	,
(	1787	)	,
(	1784	)	,
(	1781	)	,
(	1778	)	,
(	1775	)	,
(	1772	)	,
(	1769	)	,
(	1767	)	,
(	1764	)	,
(	1761	)	,
(	1758	)	,
(	1755	)	,
(	1752	)	,
(	1750	)	,
(	1747	)	,
(	1744	)	,
(	1741	)	,
(	1739	)	,
(	1736	)	,
(	1733	)	,
(	1730	)	,
(	1728	)	,
(	1725	)	,
(	1722	)	,
(	1719	)	,
(	1717	)	,
(	1714	)	,
(	1711	)	,
(	1708	)	,
(	1706	)	,
(	1703	)	,
(	1700	)	,
(	1698	)	,
(	1695	)	,
(	1692	)	,
(	1690	)	,
(	1687	)	,
(	1684	)	,
(	1682	)	,
(	1679	)	,
(	1677	)	,
(	1674	)	,
(	1671	)	,
(	1669	)	,
(	1666	)	,
(	1664	)	,
(	1661	)	,
(	1658	)	,
(	1656	)	,
(	1653	)	,
(	1651	)	,
(	1648	)	,
(	1646	)	,
(	1643	)	,
(	1641	)	,
(	1638	)	,
(	1636	)	,
(	1633	)	,
(	1631	)	,
(	1628	)	,
(	1626	)	,
(	1623	)	,
(	1621	)	,
(	1618	)	,
(	1616	)	,
(	1613	)	,
(	1611	)	,
(	1608	)	,
(	1606	)	,
(	1603	)	,
(	1601	)	,
(	1599	)	,
(	1596	)	,
(	1594	)	,
(	1591	)	,
(	1589	)	,
(	1586	)	,
(	1584	)	,
(	1582	)	,
(	1579	)	,
(	1577	)	,
(	1575	)	,
(	1572	)	,
(	1570	)	,
(	1568	)	,
(	1565	)	,
(	1563	)	,
(	1561	)	,
(	1558	)	,
(	1556	)	,
(	1554	)	,
(	1551	)	,
(	1549	)	,
(	1547	)	,
(	1544	)	,
(	1542	)	,
(	1540	)	,
(	1538	)	,
(	1535	)	,
(	1533	)	,
(	1531	)	,
(	1528	)	,
(	1526	)	,
(	1524	)	,
(	1522	)	,
(	1520	)	,
(	1517	)	,
(	1515	)	,
(	1513	)	,
(	1511	)	,
(	1509	)	,
(	1506	)	,
(	1504	)	,
(	1502	)	,
(	1500	)	,
(	1498	)	,
(	1495	)	,
(	1493	)	,
(	1491	)	,
(	1489	)	,
(	1487	)	,
(	1485	)	,
(	1483	)	,
(	1480	)	,
(	1478	)	,
(	1476	)	,
(	1474	)	,
(	1472	)	,
(	1470	)	,
(	1468	)	,
(	1466	)	,
(	1464	)	,
(	1462	)	,
(	1459	)	,
(	1457	)	,
(	1455	)	,
(	1453	)	,
(	1451	)	,
(	1449	)	,
(	1447	)	,
(	1445	)	,
(	1443	)	,
(	1441	)	,
(	1439	)	,
(	1437	)	,
(	1435	)	,
(	1433	)	,
(	1431	)	,
(	1429	)	,
(	1427	)	,
(	1425	)	,
(	1423	)	,
(	1421	)	,
(	1419	)	,
(	1417	)	,
(	1415	)	,
(	1413	)	,
(	1411	)	,
(	1409	)	,
(	1408	)	,
(	1406	)	,
(	1404	)	,
(	1402	)	,
(	1400	)	,
(	1398	)	,
(	1396	)	,
(	1394	)	,
(	1392	)	,
(	1390	)	,
(	1388	)	,
(	1387	)	,
(	1385	)	,
(	1383	)	,
(	1381	)	,
(	1379	)	,
(	1377	)	,
(	1375	)	,
(	1374	)	,
(	1372	)	,
(	1370	)	,
(	1368	)	,
(	1366	)	,
(	1364	)	,
(	1363	)	,
(	1361	)	,
(	1359	)	,
(	1357	)	,
(	1355	)	,
(	1354	)	,
(	1352	)	,
(	1350	)	,
(	1348	)	,
(	1346	)	,
(	1345	)	,
(	1343	)	,
(	1341	)	,
(	1339	)	,
(	1338	)	,
(	1336	)	,
(	1334	)	,
(	1332	)	,
(	1331	)	,
(	1329	)	,
(	1327	)	,
(	1326	)	,
(	1324	)	,
(	1322	)	,
(	1320	)	,
(	1319	)	,
(	1317	)	,
(	1315	)	,
(	1314	)	,
(	1312	)	,
(	1310	)	,
(	1309	)	,
(	1307	)	,
(	1305	)	,
(	1304	)	,
(	1302	)	,
(	1300	)	,
(	1299	)	,
(	1297	)	,
(	1295	)	,
(	1294	)	,
(	1292	)	,
(	1291	)	,
(	1289	)	,
(	1287	)	,
(	1286	)	,
(	1284	)	,
(	1283	)	,
(	1281	)	,
(	1279	)	,
(	1278	)	,
(	1276	)	,
(	1275	)	,
(	1273	)	,
(	1271	)	,
(	1270	)	,
(	1268	)	,
(	1267	)	,
(	1265	)	,
(	1264	)	,
(	1262	)	,
(	1261	)	,
(	1259	)	,
(	1257	)	,
(	1256	)	,
(	1254	)	,
(	1253	)	,
(	1251	)	,
(	1250	)	,
(	1248	)	,
(	1247	)	,
(	1245	)	,
(	1244	)	,
(	1242	)	,
(	1241	)	,
(	1239	)	,
(	1238	)	,
(	1236	)	,
(	1235	)	,
(	1234	)	,
(	1232	)	,
(	1231	)	,
(	1229	)	,
(	1228	)	,
(	1226	)	,
(	1225	)	,
(	1223	)	,
(	1222	)	,
(	1221	)	,
(	1219	)	,
(	1218	)	,
(	1216	)	,
(	1215	)	,
(	1213	)	,
(	1212	)	,
(	1211	)	,
(	1209	)	,
(	1208	)	,
(	1206	)	,
(	1205	)	,
(	1204	)	,
(	1202	)	,
(	1201	)	,
(	1200	)	,
(	1198	)	,
(	1197	)	,
(	1195	)	,
(	1194	)	,
(	1193	)	,
(	1191	)	,
(	1190	)	,
(	1189	)	,
(	1187	)	,
(	1186	)	,
(	1185	)	,
(	1183	)	,
(	1182	)	,
(	1181	)	,
(	1179	)	,
(	1178	)	,
(	1177	)	,
(	1176	)	,
(	1174	)	,
(	1173	)	,
(	1172	)	,
(	1170	)	,
(	1169	)	,
(	1168	)	,
(	1166	)	,
(	1165	)	,
(	1164	)	,
(	1163	)	,
(	1161	)	,
(	1160	)	,
(	1159	)	,
(	1158	)	,
(	1156	)	,
(	1155	)	,
(	1154	)	,
(	1153	)	,
(	1151	)	,
(	1150	)	,
(	1149	)	,
(	1148	)	,
(	1147	)	,
(	1145	)	,
(	1144	)	,
(	1143	)	,
(	1142	)	,
(	1140	)	,
(	1139	)	,
(	1138	)	,
(	1137	)	,
(	1136	)	,
(	1134	)	,
(	1133	)	,
(	1132	)	,
(	1131	)	,
(	1130	)	,
(	1129	)	,
(	1127	)	,
(	1126	)	,
(	1125	)	,
(	1124	)	,
(	1123	)	,
(	1122	)	,
(	1120	)	,
(	1119	)	,
(	1118	)	,
(	1117	)	,
(	1116	)	,
(	1115	)	,
(	1114	)	,
(	1112	)	,
(	1111	)	,
(	1110	)	,
(	1109	)	,
(	1108	)	,
(	1107	)	,
(	1106	)	,
(	1105	)	,
(	1104	)	,
(	1102	)	,
(	1101	)	,
(	1100	)	,
(	1099	)	,
(	1098	)	,
(	1097	)	,
(	1096	)	,
(	1095	)	,
(	1094	)	,
(	1093	)	,
(	1092	)	,
(	1091	)	,
(	1090	)	,
(	1088	)	,
(	1087	)	,
(	1086	)	,
(	1085	)	,
(	1084	)	,
(	1083	)	,
(	1082	)	,
(	1081	)	,
(	1080	)	,
(	1079	)	,
(	1078	)	,
(	1077	)	,
(	1076	)	,
(	1075	)	,
(	1074	)	,
(	1073	)	,
(	1072	)	,
(	1071	)	,
(	1070	)	,
(	1069	)	,
(	1068	)	,
(	1067	)	,
(	1066	)	,
(	1065	)	,
(	1064	)	,
(	1063	)	,
(	1062	)	,
(	1061	)	,
(	1060	)	,
(	1059	)	,
(	1058	)	,
(	1057	)	,
(	1056	)	,
(	1055	)	,
(	1054	)	,
(	1053	)	,
(	1052	)	,
(	1051	)	,
(	1050	)	,
(	1049	)	,
(	1048	)	,
(	1047	)	,
(	1047	)	,
(	1046	)	,
(	1045	)	,
(	1044	)	,
(	1043	)	,
(	1042	)	,
(	1041	)	,
(	1040	)	,
(	1039	)	,
(	1038	)	,
(	1037	)	,
(	1036	)	,
(	1035	)	,
(	1035	)	,
(	1034	)	,
(	1033	)	,
(	1032	)	,
(	1031	)	,
(	1030	)	,
(	1029	)	,
(	1028	)	,
(	1027	)	,
(	1026	)	,
(	1026	)	,
(	1025	)	,
(	1024	)	,
(	1023	)	,
(	1022	)	,
(	1021	)	,
(	1020	)	,
(	1019	)	,
(	1019	)	,
(	1018	)	,
(	1017	)	,
(	1016	)	,
(	1015	)	,
(	1014	)	,
(	1014	)	,
(	1013	)	,
(	1012	)	,
(	1011	)	,
(	1010	)	,
(	1009	)	,
(	1008	)	,
(	1008	)	,
(	1007	)	,
(	1006	)	,
(	1005	)	,
(	1004	)	,
(	1003	)	,
(	1003	)	,
(	1002	)	,
(	1001	)	,
(	1000	)	,
(	999	)	,
(	999	)	,
(	998	)	,
(	997	)	,
(	996	)	,
(	995	)	,
(	995	)	,
(	994	)	,
(	993	)	,
(	992	)	,
(	991	)	,
(	991	)	,
(	990	)	,
(	989	)	,
(	988	)	,
(	988	)	,
(	987	)	,
(	986	)	,
(	985	)	,
(	984	)	,
(	984	)	,
(	983	)	,
(	982	)	,
(	981	)	,
(	981	)	,
(	980	)	,
(	979	)	,
(	978	)	,
(	978	)	,
(	977	)	,
(	976	)	,
(	975	)	,
(	975	)	,
(	974	)	,
(	973	)	,
(	972	)	,
(	972	)	,
(	971	)	,
(	970	)	,
(	969	)	,
(	969	)	,
(	968	)	,
(	967	)	,
(	967	)	,
(	966	)	,
(	965	)	,
(	964	)	,
(	964	)	,
(	963	)	,
(	962	)	,
(	962	)	,
(	961	)	,
(	960	)	,
(	959	)	,
(	959	)	,
(	958	)	,
(	957	)	,
(	957	)	,
(	956	)	,
(	955	)	,
(	955	)	,
(	954	)	,
(	953	)	,
(	953	)	,
(	952	)	,
(	951	)	,
(	950	)	,
(	950	)	,
(	949	)	,
(	948	)	,
(	948	)	,
(	947	)	,
(	946	)	,
(	946	)	,
(	945	)	,
(	944	)	,
(	944	)	,
(	943	)	,
(	942	)	,
(	942	)	,
(	941	)	,
(	941	)	,
(	940	)	,
(	939	)	,
(	939	)	,
(	938	)	,
(	937	)	,
(	937	)	,
(	936	)	,
(	935	)	,
(	935	)	,
(	934	)	,
(	933	)	,
(	933	)	,
(	932	)	,
(	932	)	,
(	931	)	,
(	930	)	,
(	930	)	,
(	929	)	,
(	928	)	,
(	928	)	,
(	927	)	,
(	927	)	,
(	926	)	,
(	925	)	,
(	925	)	,
(	924	)	,
(	923	)	,
(	923	)	,
(	922	)	,
(	922	)	,
(	921	)	,
(	920	)	,
(	920	)	,
(	919	)	,
(	919	)	,
(	918	)	,
(	917	)	,
(	917	)	,
(	916	)	,
(	916	)	,
(	915	)	,
(	914	)	,
(	914	)	,
(	913	)	,
(	913	)	,
(	912	)	,
(	912	)	,
(	911	)	,
(	910	)	,
(	910	)	,
(	909	)	,
(	909	)	,
(	908	)	,
(	908	)	,
(	907	)	,
(	906	)	,
(	906	)	,
(	905	)	,
(	905	)	,
(	904	)	,
(	904	)	,
(	903	)	,
(	902	)	,
(	902	)	,
(	901	)	,
(	901	)	,
(	900	)	,
(	900	)	,
(	899	)	,
(	899	)	,
(	898	)	,
(	897	)	,
(	897	)	,
(	896	)	,
(	896	)	,
(	895	)	,
(	895	)	,
(	894	)	,
(	894	)	,
(	893	)	,
(	893	)	,
(	892	)	,
(	891	)	,
(	891	)	,
(	890	)	,
(	890	)	,
(	889	)	,
(	889	)	,
(	888	)	,
(	888	)	,
(	887	)	,
(	887	)	,
(	886	)	,
(	886	)	,
(	885	)	,
(	885	)	,
(	884	)	,
(	884	)	,
(	883	)	,
(	882	)	,
(	882	)	,
(	881	)	,
(	881	)	,
(	880	)	,
(	880	)	,
(	879	)	,
(	879	)	,
(	878	)	,
(	878	)	,
(	877	)	,
(	877	)	,
(	876	)	,
(	876	)	,
(	875	)	,
(	875	)	,
(	874	)	,
(	874	)	,
(	873	)	,
(	873	)	,
(	872	)	,
(	872	)	,
(	871	)	,
(	871	)	,
(	870	)	,
(	870	)	,
(	869	)	,
(	869	)	,
(	868	)	,
(	868	)	,
(	867	)	,
(	867	)	,
(	866	)	,
(	866	)	,
(	865	)	,
(	865	)	,
(	865	)	,
(	864	)	,
(	864	)	,
(	863	)	,
(	863	)	,
(	862	)	,
(	862	)	,
(	861	)	,
(	861	)	,
(	860	)	,
(	860	)	,
(	859	)	,
(	859	)	,
(	858	)	,
(	858	)	,
(	857	)	,
(	857	)	,
(	856	)	,
(	856	)	,
(	855	)	,
(	855	)	,
(	855	)	,
(	854	)	,
(	854	)	,
(	853	)	,
(	853	)	,
(	852	)	,
(	852	)	,
(	851	)	,
(	851	)	,
(	850	)	,
(	850	)	,
(	849	)	,
(	849	)	,
(	849	)	,
(	848	)	,
(	848	)	,
(	847	)	,
(	847	)	,
(	846	)	,
(	846	)	,
(	845	)	,
(	845	)	,
(	844	)	,
(	844	)	,
(	844	)	,
(	843	)	,
(	843	)	,
(	842	)	,
(	842	)	,
(	841	)	,
(	841	)	,
(	840	)	,
(	840	)	,
(	840	)	,
(	839	)	,
(	839	)	,
(	838	)	,
(	838	)	,
(	837	)	,
(	837	)	,
(	836	)	,
(	836	)	,
(	836	)	,
(	835	)	,
(	835	)	,
(	834	)	,
(	834	)	,
(	833	)	,
(	833	)	,
(	833	)	,
(	832	)	,
(	832	)	,
(	831	)	,
(	831	)	,
(	830	)	,
(	830	)	,
(	830	)	,
(	829	)	,
(	829	)	,
(	828	)	,
(	828	)	,
(	827	)	,
(	827	)	,
(	827	)	,
(	826	)	,
(	826	)	,
(	825	)	,
(	825	)	,
(	824	)	,
(	824	)	,
(	824	)	,
(	823	)	,
(	823	)	,
(	822	)	,
(	822	)	,
(	821	)	,
(	821	)	,
(	821	)	,
(	820	)	,
(	820	)	,
(	819	)	,
(	819	)	,
(	819	)	,
(	818	)	,
(	818	)	,
(	817	)	,
(	817	)	,
(	816	)	,
(	816	)	,
(	816	)	,
(	815	)	,
(	815	)	,
(	814	)	,
(	814	)	,
(	814	)	,
(	813	)	,
(	813	)	,
(	812	)	,
(	812	)	,
(	812	)	,
(	811	)	,
(	811	)	,
(	810	)	,
(	810	)	,
(	809	)	,
(	809	)	,
(	809	)	,
(	808	)	,
(	808	)	,
(	807	)	,
(	807	)	,
(	807	)	,
(	806	)	,
(	806	)	,
(	805	)	,
(	805	)	,
(	805	)	,
(	804	)	,
(	804	)	,
(	803	)	,
(	803	)	,
(	803	)	,
(	802	)	,
(	802	)	,
(	801	)	,
(	801	)	,
(	801	)	,
(	800	)	,
(	800	)	,
(	799	)	,
(	799	)	,
(	799	)	,
(	798	)	,
(	798	)	,
(	797	)	,
(	797	)	,
(	797	)	,
(	796	)	,
(	796	)	,
(	795	)	,
(	795	)	,
(	795	)	,
(	794	)	,
(	794	)	,
(	793	)	,
(	793	)	,
(	793	)	,
(	792	)	,
(	792	)	,
(	791	)	,
(	791	)	,
(	791	)	,
(	790	)	,
(	790	)	,
(	789	)	,
(	789	)	,
(	789	)	,
(	788	)	,
(	788	)	,
(	787	)	,
(	787	)	,
(	787	)	,
(	786	)	,
(	786	)	,
(	785	)	,
(	785	)	,
(	785	)	,
(	784	)	,
(	784	)	,
(	783	)	,
(	783	)	,
(	783	)	,
(	782	)	,
(	782	)	,
(	781	)	,
(	781	)	,
(	781	)	,
(	780	)	,
(	780	)	,
(	779	)	,
(	779	)	,
(	779	)	,
(	778	)	,
(	778	)	,
(	777	)	,
(	777	)	,
(	777	)	,
(	776	)	,
(	776	)	,
(	776	)	,
(	775	)	,
(	775	)	,
(	774	)	,
(	774	)	,
(	774	)	,
(	773	)	,
(	773	)	,
(	772	)	,
(	772	)	,
(	772	)	,
(	771	)	,
(	771	)	,
(	770	)	,
(	770	)	,
(	770	)	,
(	769	)	,
(	769	)	,
(	768	)	,
(	768	)	,
(	768	)	,
(	767	)	,
(	767	)	,
(	766	)	,
(	766	)	,
(	766	)	,
(	765	)	,
(	765	)	,
(	764	)	,
(	764	)	,
(	764	)	,
(	763	)	,
(	763	)	,
(	763	)	,
(	762	)	,
(	762	)	,
(	761	)	,
(	761	)	,
(	761	)	,
(	760	)	,
(	760	)	,
(	759	)	,
(	759	)	,
(	759	)	,
(	758	)	,
(	758	)	,
(	757	)	,
(	757	)	,
(	757	)	,
(	756	)	,
(	756	)	,
(	755	)	,
(	755	)	,
(	755	)	,
(	754	)	,
(	754	)	,
(	753	)	,
(	753	)	,
(	753	)	,
(	752	)	,
(	752	)	,
(	752	)	,
(	751	)	,
(	751	)	,
(	750	)	,
(	750	)	,
(	750	)	,
(	749	)	,
(	749	)	,
(	748	)	,
(	748	)	,
(	748	)	,
(	747	)	,
(	747	)	,
(	746	)	,
(	746	)	,
(	746	)	,
(	745	)	,
(	745	)	,
(	744	)	,
(	744	)	,
(	744	)	,
(	743	)	,
(	743	)	,
(	742	)	,
(	742	)	,
(	742	)	,
(	741	)	,
(	741	)	,
(	740	)	,
(	740	)	,
(	740	)	,
(	739	)	,
(	739	)	,
(	738	)	,
(	738	)	,
(	738	)	,
(	737	)	,
(	737	)	,
(	736	)	,
(	736	)	,
(	736	)	,
(	735	)	,
(	735	)	,
(	734	)	,
(	734	)	,
(	734	)	,
(	733	)	,
(	733	)	,
(	732	)	,
(	732	)	,
(	732	)	,
(	731	)	,
(	731	)	,
(	730	)	,
(	730	)	,
(	730	)	,
(	729	)	,
(	729	)	,
(	728	)	,
(	728	)	,
(	728	)	,
(	727	)	,
(	727	)	,
(	726	)	,
(	726	)	,
(	726	)	,
(	725	)	,
(	725	)	,
(	724	)	,
(	724	)	,
(	724	)	,
(	723	)	,
(	723	)	,
(	722	)	,
(	722	)	,
(	722	)	,
(	721	)	,
(	721	)	,
(	720	)	,
(	720	)	,
(	720	)	,
(	719	)	,
(	719	)	,
(	718	)	,
(	718	)	,
(	717	)	,
(	717	)	,
(	717	)	,
(	716	)	,
(	716	)	,
(	715	)	,
(	715	)	,
(	715	)	,
(	714	)	,
(	714	)	,
(	713	)	,
(	713	)	,
(	713	)	,
(	712	)	,
(	712	)	,
(	711	)	,
(	711	)	,
(	710	)	,
(	710	)	,
(	710	)	,
(	709	)	,
(	709	)	,
(	708	)	,
(	708	)	,
(	708	)	,
(	707	)	,
(	707	)	,
(	706	)	,
(	706	)	,
(	706	)	,
(	705	)	,
(	705	)	,
(	704	)	,
(	704	)	,
(	703	)	,
(	703	)	,
(	703	)	,
(	702	)	,
(	702	)	,
(	701	)	,
(	701	)	,
(	701	)	,
(	700	)	,
(	700	)	,
(	699	)	,
(	699	)	,
(	698	)	,
(	698	)	,
(	698	)	,
(	697	)	,
(	697	)	,
(	696	)	,
(	696	)	,
(	695	)	,
(	695	)	,
(	695	)	,
(	694	)	,
(	694	)	,
(	693	)	,
(	693	)	,
(	693	)	,
(	692	)	,
(	692	)	,
(	691	)	,
(	691	)	,
(	690	)	,
(	690	)	,
(	690	)	,
(	689	)	,
(	689	)	,
(	688	)	,
(	688	)	,
(	687	)	,
(	687	)	,
(	687	)	,
(	686	)	,
(	686	)	,
(	685	)	,
(	685	)	,
(	684	)	,
(	684	)	,
(	684	)	,
(	683	)	,
(	683	)	,
(	682	)	,
(	682	)	,
(	681	)	,
(	681	)	,
(	681	)	,
(	680	)	,
(	680	)	,
(	679	)	,
(	679	)	,
(	678	)	,
(	678	)	,
(	678	)	,
(	677	)	,
(	677	)	,
(	676	)	,
(	676	)	,
(	675	)	,
(	675	)	,
(	674	)	,
(	674	)	,
(	674	)	,
(	673	)	,
(	673	)	,
(	672	)	,
(	672	)	,
(	671	)	,
(	671	)	,
(	671	)	,
(	670	)	,
(	670	)	,
(	669	)	,
(	669	)	,
(	668	)	,
(	668	)	,
(	667	)	,
(	667	)	,
(	667	)	,
(	666	)	,
(	666	)	,
(	665	)	,
(	665	)	,
(	664	)	,
(	664	)	,
(	664	)	,
(	663	)	,
(	663	)	,
(	662	)	,
(	662	)	,
(	661	)	,
(	661	)	,
(	660	)	,
(	660	)	,
(	660	)	,
(	659	)	,
(	659	)	,
(	658	)	,
(	658	)	,
(	657	)	,
(	657	)	,
(	656	)	,
(	656	)	,
(	655	)	,
(	655	)	,
(	655	)	,
(	654	)	,
(	654	)	,
(	653	)	,
(	653	)	,
(	652	)	,
(	652	)	,
(	651	)	,
(	651	)	,
(	651	)	,
(	650	)	,
(	650	)	,
(	649	)	,
(	649	)	,
(	648	)	,
(	648	)	,
(	647	)	,
(	647	)	,
(	646	)	,
(	646	)	,
(	646	)	,
(	645	)	,
(	645	)	,
(	644	)	,
(	644	)	,
(	643	)	,
(	643	)	,
(	642	)	,
(	642	)	,
(	641	)	,
(	641	)	,
(	641	)	,
(	640	)	,
(	640	)	,
(	639	)	,
(	639	)	,
(	638	)	,
(	638	)	,
(	637	)	,
(	637	)	,
(	636	)	,
(	636	)	,
(	636	)	,
(	635	)	,
(	635	)	,
(	634	)	,
(	634	)	,
(	633	)	,
(	633	)	,
(	632	)	,
(	632	)	,
(	631	)	,
(	631	)	,
(	630	)	,
(	630	)	,
(	630	)	,
(	629	)	,
(	629	)	,
(	628	)	,
(	628	)	,
(	627	)	,
(	627	)	,
(	626	)	,
(	626	)	,
(	625	)	,
(	625	)	,
(	624	)	,
(	624	)	,
(	624	)	,
(	623	)	,
(	623	)	,
(	622	)	,
(	622	)	,
(	621	)	,
(	621	)	,
(	620	)	,
(	620	)	,
(	619	)	,
(	619	)	,
(	618	)	,
(	618	)	,
(	617	)	,
(	617	)	,
(	616	)	,
(	616	)	,
(	616	)	,
(	615	)	,
(	615	)	,
(	614	)	,
(	614	)	,
(	613	)	,
(	613	)	,
(	612	)	,
(	612	)	,
(	611	)	,
(	611	)	,
(	610	)	,
(	610	)	,
(	609	)	,
(	609	)	,
(	609	)	,
(	608	)	,
(	608	)	,
(	607	)	,
(	607	)	,
(	606	)	,
(	606	)	,
(	605	)	,
(	605	)	,
(	604	)	,
(	604	)	,
(	603	)	,
(	603	)	,
(	602	)	,
(	602	)	,
(	601	)	,
(	601	)	,
(	600	)	,
(	600	)	,
(	600	)	,
(	599	)	,
(	599	)	,
(	598	)	,
(	598	)	,
(	597	)	,
(	597	)	,
(	596	)	,
(	596	)	,
(	595	)	,
(	595	)	,
(	594	)	,
(	594	)	,
(	593	)	,
(	593	)	,
(	592	)	,
(	592	)	,
(	591	)	,
(	591	)	,
(	590	)	,
(	590	)	,
(	590	)	,
(	589	)	,
(	589	)	,
(	588	)	,
(	588	)	,
(	587	)	,
(	587	)	,
(	586	)	,
(	586	)	,
(	585	)	,
(	585	)	,
(	584	)	,
(	584	)	,
(	583	)	,
(	583	)	,
(	582	)	,
(	582	)	,
(	581	)	,
(	581	)	,
(	580	)	,
(	580	)	,
(	579	)	,
(	579	)	,
(	578	)	,
(	578	)	,
(	578	)	,
(	577	)	,
(	577	)	,
(	576	)	,
(	576	)	,
(	575	)	,
(	575	)	,
(	574	)	,
(	574	)	,
(	573	)	,
(	573	)	,
(	572	)	,
(	572	)	,
(	571	)	,
(	571	)	,
(	570	)	,
(	570	)	,
(	569	)	,
(	569	)	,
(	568	)	,
(	568	)	,
(	567	)	,
(	567	)	,
(	566	)	,
(	566	)	,
(	566	)	,
(	565	)	,
(	565	)	,
(	564	)	,
(	564	)	,
(	563	)	,
(	563	)	,
(	562	)	,
(	562	)	,
(	561	)	,
(	561	)	,
(	560	)	,
(	560	)	,
(	559	)	,
(	559	)	,
(	558	)	,
(	558	)	,
(	557	)	,
(	557	)	,
(	556	)	,
(	556	)	,
(	555	)	,
(	555	)	,
(	554	)	,
(	554	)	,
(	554	)	,
(	553	)	,
(	553	)	,
(	552	)	,
(	552	)	,
(	551	)	,
(	551	)	,
(	550	)	,
(	550	)	,
(	549	)	,
(	549	)	,
(	548	)	,
(	548	)	,
(	547	)	,
(	547	)	,
(	546	)	,
(	546	)	,
(	545	)	,
(	545	)	,
(	544	)	,
(	544	)	,
(	543	)	,
(	543	)	,
(	543	)	,
(	542	)	,
(	542	)	,
(	541	)	,
(	541	)	,
(	540	)	,
(	540	)	,
(	539	)	,
(	539	)	,
(	538	)	,
(	538	)	,
(	537	)	,
(	537	)	,
(	536	)	,
(	536	)	,
(	535	)	,
(	535	)	,
(	534	)	,
(	534	)	,
(	534	)	,
(	533	)	,
(	533	)	,
(	532	)	,
(	532	)	,
(	531	)	,
(	531	)	,
(	530	)	,
(	530	)	,
(	529	)	,
(	529	)	,
(	528	)	,
(	528	)	,
(	527	)	,
(	527	)	,
(	526	)	,
(	526	)	,
(	525	)	,
(	525	)	,
(	525	)	,
(	524	)	,
(	524	)	,
(	523	)	,
(	523	)	,
(	522	)	,
(	522	)	,
(	521	)	,
(	521	)	,
(	520	)	,
(	520	)	,
(	519	)	,
(	519	)	,
(	518	)	,
(	518	)	,
(	518	)	,
(	517	)	,
(	517	)	,
(	516	)	,
(	516	)	,
(	515	)	,
(	515	)	,
(	514	)	,
(	514	)	,
(	513	)	,
(	513	)	,
(	512	)	,
(	512	)	,
(	512	)	,
(	511	)	,
(	511	)	,
(	510	)	,
(	510	)	,
(	509	)	,
(	509	)	,
(	508	)	,
(	508	)	,
(	507	)	,
(	507	)	,
(	506	)	,
(	506	)	,
(	506	)	,
(	505	)	,
(	505	)	,
(	504	)	,
(	504	)	,
(	503	)	,
(	503	)	,
(	502	)	,
(	502	)	,
(	501	)	,
(	501	)	,
(	501	)	,
(	500	)	,
(	500	)	,
(	499	)	,
(	499	)	,
(	498	)	,
(	498	)	,
(	497	)	,
(	497	)	,
(	497	)	,
(	496	)	,
(	496	)	,
(	495	)	,
(	495	)	,
(	494	)	,
(	494	)	,
(	493	)	,
(	493	)	,
(	493	)	,
(	492	)	,
(	492	)	,
(	491	)	,
(	491	)	,
(	490	)	,
(	490	)	,
(	489	)	,
(	489	)	,
(	489	)	,
(	488	)	,
(	488	)	,
(	487	)	,
(	487	)	,
(	486	)	,
(	486	)	,
(	486	)	,
(	485	)	,
(	485	)	,
(	484	)	,
(	484	)	,
(	483	)	,
(	483	)	,
(	483	)	,
(	482	)	,
(	482	)	,
(	481	)	,
(	481	)	,
(	480	)	,
(	480	)	,
(	480	)	,
(	479	)	,
(	479	)	,
(	478	)	,
(	478	)	,
(	477	)	,
(	477	)	,
(	477	)	,
(	476	)	,
(	476	)	,
(	475	)	,
(	475	)	,
(	475	)	,
(	474	)	,
(	474	)	,
(	473	)	,
(	473	)	,
(	472	)	,
(	472	)	,
(	472	)	,
(	471	)	,
(	471	)	,
(	470	)	,
(	470	)	,
(	470	)	,
(	469	)	,
(	469	)	,
(	468	)	,
(	468	)	,
(	468	)	,
(	467	)	,
(	467	)	,
(	466	)	,
(	466	)	,
(	466	)	,
(	465	)	,
(	465	)	,
(	464	)	,
(	464	)	,
(	464	)	,
(	463	)	,
(	463	)	,
(	462	)	,
(	462	)	,
(	462	)	,
(	461	)	,
(	461	)	,
(	460	)	,
(	460	)	,
(	460	)	,
(	459	)	,
(	459	)	,
(	459	)	,
(	458	)	,
(	458	)	,
(	457	)	,
(	457	)	,
(	457	)	,
(	456	)	,
(	456	)	,
(	455	)	,
(	455	)	,
(	455	)	,
(	454	)	,
(	454	)	,
(	454	)	,
(	453	)	,
(	453	)	,
(	453	)	,
(	452	)	,
(	452	)	,
(	451	)	,
(	451	)	,
(	451	)	,
(	450	)	,
(	450	)	,
(	450	)	,
(	449	)	,
(	449	)	,
(	449	)	,
(	448	)	,
(	448	)	,
(	447	)	,
(	447	)	,
(	447	)	,
(	446	)	,
(	446	)	,
(	446	)	,
(	445	)	,
(	445	)	,
(	445	)	,
(	444	)	,
(	444	)	,
(	444	)	,
(	443	)	,
(	443	)	,
(	443	)	,
(	442	)	,
(	442	)	,
(	442	)	,
(	441	)	,
(	441	)	,
(	441	)	,
(	440	)	,
(	440	)	,
(	440	)	,
(	439	)	,
(	439	)	,
(	439	)	,
(	438	)	,
(	438	)	,
(	438	)	,
(	437	)	,
(	437	)	,
(	437	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	436	)	,
(	435	)	,
(	435	)	,
(	435	)	,
(	434	)	,
(	434	)	,
(	434	)	,
(	433	)	,
(	433	)	,
(	433	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	432	)	,
(	431	)	,
(	431	)	,
(	431	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	430	)	,
(	429	)	,
(	429	)	,
(	429	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	428	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	427	)	,
(	426	)	,
(	426	)	,
(	426	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	425	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	424	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	423	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	422	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	421	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	420	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	419	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	418	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	417	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	416	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	415	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	414	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	413	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	412	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	411	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	410	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	409	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	408	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	407	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	406	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	405	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	404	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	403	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	402	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	401	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	,
(	400	)	





);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
    	
   distance <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),distance'length));
	
end behavior;

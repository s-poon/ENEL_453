
-- In this example, we're going to map voltage to distance, using a linear 
-- approximation, according to the Sharp GP2Y0A41SK0F datasheet page 4, or 
-- Lab 3 handout page 5. 
-- 
-- The relevant points we will select are:
-- 2.750 V is  4.00 cm (or 2750 mV and  40.0 mm)
-- 0.400 V is 33.00 cm (or  400 mV and 330.0 mm)
-- 
-- Mapping to the scales in our system
-- 2750 (mV) should map to  400 (10^-4 m)
--  400 (mV) should map to 3300 (10^-4 m)
-- and developing a linear equation, we find:
--
-- Distance = -2900/2350 * Voltage + 3793.617
-- Note this code implements linear function, you must map to the 
-- NON-linear relationship in the datasheet. This code is only provided 
-- for reference to help get you started.

LIBRARY ieee;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

ENTITY dis2freq IS
   PORT(
      clk            :  IN    STD_LOGIC;                                
      reset          :  IN    STD_LOGIC;                                
      voltage        :  IN    STD_LOGIC_VECTOR(12 DOWNTO 0);                           
      frequency       :  OUT   STD_LOGIC_VECTOR(14 DOWNTO 0));  
END dis2freq;

ARCHITECTURE behavior OF dis2freq IS

-- This array has been pasted in from the Excel spreadsheet.
-- In this array, the values are distances, in units 10^-4 m. 
-- To get cm, move the decimal point 2 places to the left.
-- See how to get the distance output at the bottom of this file,
-- after begin.

type array_1d is array (0 to 4095) of integer;
constant v2d_LUT : array_1d := (

(	2250	)	,
(	2251	)	,
(	2251	)	,
(	2252	)	,
(	2252	)	,
(	2253	)	,
(	2253	)	,
(	2254	)	,
(	2255	)	,
(	2255	)	,
(	2256	)	,
(	2256	)	,
(	2257	)	,
(	2257	)	,
(	2258	)	,
(	2258	)	,
(	2259	)	,
(	2260	)	,
(	2260	)	,
(	2261	)	,
(	2261	)	,
(	2262	)	,
(	2262	)	,
(	2263	)	,
(	2264	)	,
(	2264	)	,
(	2265	)	,
(	2265	)	,
(	2266	)	,
(	2266	)	,
(	2267	)	,
(	2268	)	,
(	2268	)	,
(	2269	)	,
(	2269	)	,
(	2270	)	,
(	2270	)	,
(	2271	)	,
(	2272	)	,
(	2272	)	,
(	2273	)	,
(	2273	)	,
(	2274	)	,
(	2274	)	,
(	2275	)	,
(	2276	)	,
(	2276	)	,
(	2277	)	,
(	2277	)	,
(	2278	)	,
(	2278	)	,
(	2279	)	,
(	2280	)	,
(	2280	)	,
(	2281	)	,
(	2281	)	,
(	2282	)	,
(	2283	)	,
(	2283	)	,
(	2284	)	,
(	2284	)	,
(	2285	)	,
(	2285	)	,
(	2286	)	,
(	2287	)	,
(	2287	)	,
(	2288	)	,
(	2288	)	,
(	2289	)	,
(	2289	)	,
(	2290	)	,
(	2291	)	,
(	2291	)	,
(	2292	)	,
(	2292	)	,
(	2293	)	,
(	2294	)	,
(	2294	)	,
(	2295	)	,
(	2295	)	,
(	2296	)	,
(	2297	)	,
(	2297	)	,
(	2298	)	,
(	2298	)	,
(	2299	)	,
(	2299	)	,
(	2300	)	,
(	2301	)	,
(	2301	)	,
(	2302	)	,
(	2302	)	,
(	2303	)	,
(	2304	)	,
(	2304	)	,
(	2305	)	,
(	2305	)	,
(	2306	)	,
(	2307	)	,
(	2307	)	,
(	2308	)	,
(	2308	)	,
(	2309	)	,
(	2309	)	,
(	2310	)	,
(	2311	)	,
(	2311	)	,
(	2312	)	,
(	2312	)	,
(	2313	)	,
(	2314	)	,
(	2314	)	,
(	2315	)	,
(	2315	)	,
(	2316	)	,
(	2317	)	,
(	2317	)	,
(	2318	)	,
(	2318	)	,
(	2319	)	,
(	2320	)	,
(	2320	)	,
(	2321	)	,
(	2321	)	,
(	2322	)	,
(	2323	)	,
(	2323	)	,
(	2324	)	,
(	2324	)	,
(	2325	)	,
(	2326	)	,
(	2326	)	,
(	2327	)	,
(	2327	)	,
(	2328	)	,
(	2329	)	,
(	2329	)	,
(	2330	)	,
(	2330	)	,
(	2331	)	,
(	2332	)	,
(	2332	)	,
(	2333	)	,
(	2333	)	,
(	2334	)	,
(	2335	)	,
(	2335	)	,
(	2336	)	,
(	2336	)	,
(	2337	)	,
(	2338	)	,
(	2338	)	,
(	2339	)	,
(	2339	)	,
(	2340	)	,
(	2341	)	,
(	2341	)	,
(	2342	)	,
(	2343	)	,
(	2343	)	,
(	2344	)	,
(	2344	)	,
(	2345	)	,
(	2346	)	,
(	2346	)	,
(	2347	)	,
(	2347	)	,
(	2348	)	,
(	2349	)	,
(	2349	)	,
(	2350	)	,
(	2350	)	,
(	2351	)	,
(	2352	)	,
(	2352	)	,
(	2353	)	,
(	2354	)	,
(	2354	)	,
(	2355	)	,
(	2355	)	,
(	2356	)	,
(	2357	)	,
(	2357	)	,
(	2358	)	,
(	2358	)	,
(	2359	)	,
(	2360	)	,
(	2360	)	,
(	2361	)	,
(	2362	)	,
(	2362	)	,
(	2363	)	,
(	2363	)	,
(	2364	)	,
(	2365	)	,
(	2365	)	,
(	2366	)	,
(	2367	)	,
(	2367	)	,
(	2368	)	,
(	2368	)	,
(	2369	)	,
(	2370	)	,
(	2370	)	,
(	2371	)	,
(	2372	)	,
(	2372	)	,
(	2373	)	,
(	2373	)	,
(	2374	)	,
(	2375	)	,
(	2375	)	,
(	2376	)	,
(	2377	)	,
(	2377	)	,
(	2378	)	,
(	2378	)	,
(	2379	)	,
(	2380	)	,
(	2380	)	,
(	2381	)	,
(	2382	)	,
(	2382	)	,
(	2383	)	,
(	2383	)	,
(	2384	)	,
(	2385	)	,
(	2385	)	,
(	2386	)	,
(	2387	)	,
(	2387	)	,
(	2388	)	,
(	2389	)	,
(	2389	)	,
(	2390	)	,
(	2390	)	,
(	2391	)	,
(	2392	)	,
(	2392	)	,
(	2393	)	,
(	2394	)	,
(	2394	)	,
(	2395	)	,
(	2396	)	,
(	2396	)	,
(	2397	)	,
(	2397	)	,
(	2398	)	,
(	2399	)	,
(	2399	)	,
(	2400	)	,
(	2401	)	,
(	2401	)	,
(	2402	)	,
(	2403	)	,
(	2403	)	,
(	2404	)	,
(	2404	)	,
(	2405	)	,
(	2406	)	,
(	2406	)	,
(	2407	)	,
(	2408	)	,
(	2408	)	,
(	2409	)	,
(	2410	)	,
(	2410	)	,
(	2411	)	,
(	2412	)	,
(	2412	)	,
(	2413	)	,
(	2414	)	,
(	2414	)	,
(	2415	)	,
(	2415	)	,
(	2416	)	,
(	2417	)	,
(	2417	)	,
(	2418	)	,
(	2419	)	,
(	2419	)	,
(	2420	)	,
(	2421	)	,
(	2421	)	,
(	2422	)	,
(	2423	)	,
(	2423	)	,
(	2424	)	,
(	2425	)	,
(	2425	)	,
(	2426	)	,
(	2427	)	,
(	2427	)	,
(	2428	)	,
(	2428	)	,
(	2429	)	,
(	2430	)	,
(	2430	)	,
(	2431	)	,
(	2432	)	,
(	2432	)	,
(	2433	)	,
(	2434	)	,
(	2434	)	,
(	2435	)	,
(	2436	)	,
(	2436	)	,
(	2437	)	,
(	2438	)	,
(	2438	)	,
(	2439	)	,
(	2440	)	,
(	2440	)	,
(	2441	)	,
(	2442	)	,
(	2442	)	,
(	2443	)	,
(	2444	)	,
(	2444	)	,
(	2445	)	,
(	2446	)	,
(	2446	)	,
(	2447	)	,
(	2448	)	,
(	2448	)	,
(	2449	)	,
(	2450	)	,
(	2450	)	,
(	2451	)	,
(	2452	)	,
(	2452	)	,
(	2453	)	,
(	2454	)	,
(	2454	)	,
(	2455	)	,
(	2456	)	,
(	2456	)	,
(	2457	)	,
(	2458	)	,
(	2458	)	,
(	2459	)	,
(	2460	)	,
(	2460	)	,
(	2461	)	,
(	2462	)	,
(	2462	)	,
(	2463	)	,
(	2464	)	,
(	2464	)	,
(	2465	)	,
(	2466	)	,
(	2466	)	,
(	2467	)	,
(	2468	)	,
(	2468	)	,
(	2469	)	,
(	2470	)	,
(	2470	)	,
(	2471	)	,
(	2472	)	,
(	2473	)	,
(	2473	)	,
(	2474	)	,
(	2475	)	,
(	2475	)	,
(	2476	)	,
(	2477	)	,
(	2477	)	,
(	2478	)	,
(	2479	)	,
(	2479	)	,
(	2480	)	,
(	2481	)	,
(	2481	)	,
(	2482	)	,
(	2483	)	,
(	2483	)	,
(	2484	)	,
(	2485	)	,
(	2486	)	,
(	2486	)	,
(	2487	)	,
(	2488	)	,
(	2488	)	,
(	2489	)	,
(	2490	)	,
(	2490	)	,
(	2491	)	,
(	2492	)	,
(	2492	)	,
(	2493	)	,
(	2494	)	,
(	2494	)	,
(	2495	)	,
(	2496	)	,
(	2497	)	,
(	2497	)	,
(	2498	)	,
(	2499	)	,
(	2499	)	,
(	2500	)	,
(	2501	)	,
(	2501	)	,
(	2502	)	,
(	2503	)	,
(	2503	)	,
(	2504	)	,
(	2505	)	,
(	2506	)	,
(	2506	)	,
(	2507	)	,
(	2508	)	,
(	2508	)	,
(	2509	)	,
(	2510	)	,
(	2510	)	,
(	2511	)	,
(	2512	)	,
(	2513	)	,
(	2513	)	,
(	2514	)	,
(	2515	)	,
(	2515	)	,
(	2516	)	,
(	2517	)	,
(	2517	)	,
(	2518	)	,
(	2519	)	,
(	2520	)	,
(	2520	)	,
(	2521	)	,
(	2522	)	,
(	2522	)	,
(	2523	)	,
(	2524	)	,
(	2525	)	,
(	2525	)	,
(	2526	)	,
(	2527	)	,
(	2527	)	,
(	2528	)	,
(	2529	)	,
(	2530	)	,
(	2530	)	,
(	2531	)	,
(	2532	)	,
(	2532	)	,
(	2533	)	,
(	2534	)	,
(	2534	)	,
(	2535	)	,
(	2536	)	,
(	2537	)	,
(	2537	)	,
(	2538	)	,
(	2539	)	,
(	2540	)	,
(	2540	)	,
(	2541	)	,
(	2542	)	,
(	2542	)	,
(	2543	)	,
(	2544	)	,
(	2545	)	,
(	2545	)	,
(	2546	)	,
(	2547	)	,
(	2547	)	,
(	2548	)	,
(	2549	)	,
(	2550	)	,
(	2550	)	,
(	2551	)	,
(	2552	)	,
(	2552	)	,
(	2553	)	,
(	2554	)	,
(	2555	)	,
(	2555	)	,
(	2556	)	,
(	2557	)	,
(	2558	)	,
(	2558	)	,
(	2559	)	,
(	2560	)	,
(	2560	)	,
(	2561	)	,
(	2562	)	,
(	2563	)	,
(	2563	)	,
(	2564	)	,
(	2565	)	,
(	2566	)	,
(	2566	)	,
(	2567	)	,
(	2568	)	,
(	2568	)	,
(	2569	)	,
(	2570	)	,
(	2571	)	,
(	2571	)	,
(	2572	)	,
(	2573	)	,
(	2574	)	,
(	2574	)	,
(	2575	)	,
(	2576	)	,
(	2577	)	,
(	2577	)	,
(	2578	)	,
(	2579	)	,
(	2580	)	,
(	2580	)	,
(	2581	)	,
(	2582	)	,
(	2582	)	,
(	2583	)	,
(	2584	)	,
(	2585	)	,
(	2585	)	,
(	2586	)	,
(	2587	)	,
(	2588	)	,
(	2588	)	,
(	2589	)	,
(	2590	)	,
(	2591	)	,
(	2591	)	,
(	2592	)	,
(	2593	)	,
(	2594	)	,
(	2594	)	,
(	2595	)	,
(	2596	)	,
(	2597	)	,
(	2597	)	,
(	2598	)	,
(	2599	)	,
(	2600	)	,
(	2600	)	,
(	2601	)	,
(	2602	)	,
(	2603	)	,
(	2603	)	,
(	2604	)	,
(	2605	)	,
(	2606	)	,
(	2606	)	,
(	2607	)	,
(	2608	)	,
(	2609	)	,
(	2609	)	,
(	2610	)	,
(	2611	)	,
(	2612	)	,
(	2612	)	,
(	2613	)	,
(	2614	)	,
(	2615	)	,
(	2616	)	,
(	2616	)	,
(	2617	)	,
(	2618	)	,
(	2619	)	,
(	2619	)	,
(	2620	)	,
(	2621	)	,
(	2622	)	,
(	2622	)	,
(	2623	)	,
(	2624	)	,
(	2625	)	,
(	2625	)	,
(	2626	)	,
(	2627	)	,
(	2628	)	,
(	2629	)	,
(	2629	)	,
(	2630	)	,
(	2631	)	,
(	2632	)	,
(	2632	)	,
(	2633	)	,
(	2634	)	,
(	2635	)	,
(	2635	)	,
(	2636	)	,
(	2637	)	,
(	2638	)	,
(	2639	)	,
(	2639	)	,
(	2640	)	,
(	2641	)	,
(	2642	)	,
(	2642	)	,
(	2643	)	,
(	2644	)	,
(	2645	)	,
(	2646	)	,
(	2646	)	,
(	2647	)	,
(	2648	)	,
(	2649	)	,
(	2649	)	,
(	2650	)	,
(	2651	)	,
(	2652	)	,
(	2653	)	,
(	2653	)	,
(	2654	)	,
(	2655	)	,
(	2656	)	,
(	2656	)	,
(	2657	)	,
(	2658	)	,
(	2659	)	,
(	2660	)	,
(	2660	)	,
(	2661	)	,
(	2662	)	,
(	2663	)	,
(	2664	)	,
(	2664	)	,
(	2665	)	,
(	2666	)	,
(	2667	)	,
(	2667	)	,
(	2668	)	,
(	2669	)	,
(	2670	)	,
(	2671	)	,
(	2671	)	,
(	2672	)	,
(	2673	)	,
(	2674	)	,
(	2675	)	,
(	2675	)	,
(	2676	)	,
(	2677	)	,
(	2678	)	,
(	2679	)	,
(	2679	)	,
(	2680	)	,
(	2681	)	,
(	2682	)	,
(	2683	)	,
(	2683	)	,
(	2684	)	,
(	2685	)	,
(	2686	)	,
(	2687	)	,
(	2687	)	,
(	2688	)	,
(	2689	)	,
(	2690	)	,
(	2691	)	,
(	2691	)	,
(	2692	)	,
(	2693	)	,
(	2694	)	,
(	2695	)	,
(	2695	)	,
(	2696	)	,
(	2697	)	,
(	2698	)	,
(	2699	)	,
(	2699	)	,
(	2700	)	,
(	2701	)	,
(	2702	)	,
(	2703	)	,
(	2704	)	,
(	2704	)	,
(	2705	)	,
(	2706	)	,
(	2707	)	,
(	2708	)	,
(	2708	)	,
(	2709	)	,
(	2710	)	,
(	2711	)	,
(	2712	)	,
(	2712	)	,
(	2713	)	,
(	2714	)	,
(	2715	)	,
(	2716	)	,
(	2717	)	,
(	2717	)	,
(	2718	)	,
(	2719	)	,
(	2720	)	,
(	2721	)	,
(	2721	)	,
(	2722	)	,
(	2723	)	,
(	2724	)	,
(	2725	)	,
(	2726	)	,
(	2726	)	,
(	2727	)	,
(	2728	)	,
(	2729	)	,
(	2730	)	,
(	2731	)	,
(	2731	)	,
(	2732	)	,
(	2733	)	,
(	2734	)	,
(	2735	)	,
(	2736	)	,
(	2736	)	,
(	2737	)	,
(	2738	)	,
(	2739	)	,
(	2740	)	,
(	2741	)	,
(	2741	)	,
(	2742	)	,
(	2743	)	,
(	2744	)	,
(	2745	)	,
(	2746	)	,
(	2746	)	,
(	2747	)	,
(	2748	)	,
(	2749	)	,
(	2750	)	,
(	2751	)	,
(	2751	)	,
(	2752	)	,
(	2753	)	,
(	2754	)	,
(	2755	)	,
(	2756	)	,
(	2757	)	,
(	2757	)	,
(	2758	)	,
(	2759	)	,
(	2760	)	,
(	2761	)	,
(	2762	)	,
(	2762	)	,
(	2763	)	,
(	2764	)	,
(	2765	)	,
(	2766	)	,
(	2767	)	,
(	2768	)	,
(	2768	)	,
(	2769	)	,
(	2770	)	,
(	2771	)	,
(	2772	)	,
(	2773	)	,
(	2773	)	,
(	2774	)	,
(	2775	)	,
(	2776	)	,
(	2777	)	,
(	2778	)	,
(	2779	)	,
(	2779	)	,
(	2780	)	,
(	2781	)	,
(	2782	)	,
(	2783	)	,
(	2784	)	,
(	2785	)	,
(	2786	)	,
(	2786	)	,
(	2787	)	,
(	2788	)	,
(	2789	)	,
(	2790	)	,
(	2791	)	,
(	2792	)	,
(	2792	)	,
(	2793	)	,
(	2794	)	,
(	2795	)	,
(	2796	)	,
(	2797	)	,
(	2798	)	,
(	2799	)	,
(	2799	)	,
(	2800	)	,
(	2801	)	,
(	2802	)	,
(	2803	)	,
(	2804	)	,
(	2805	)	,
(	2805	)	,
(	2806	)	,
(	2807	)	,
(	2808	)	,
(	2809	)	,
(	2810	)	,
(	2811	)	,
(	2812	)	,
(	2813	)	,
(	2813	)	,
(	2814	)	,
(	2815	)	,
(	2816	)	,
(	2817	)	,
(	2818	)	,
(	2819	)	,
(	2820	)	,
(	2820	)	,
(	2821	)	,
(	2822	)	,
(	2823	)	,
(	2824	)	,
(	2825	)	,
(	2826	)	,
(	2827	)	,
(	2828	)	,
(	2828	)	,
(	2829	)	,
(	2830	)	,
(	2831	)	,
(	2832	)	,
(	2833	)	,
(	2834	)	,
(	2835	)	,
(	2836	)	,
(	2836	)	,
(	2837	)	,
(	2838	)	,
(	2839	)	,
(	2840	)	,
(	2841	)	,
(	2842	)	,
(	2843	)	,
(	2844	)	,
(	2845	)	,
(	2845	)	,
(	2846	)	,
(	2847	)	,
(	2848	)	,
(	2849	)	,
(	2850	)	,
(	2851	)	,
(	2852	)	,
(	2853	)	,
(	2854	)	,
(	2854	)	,
(	2855	)	,
(	2856	)	,
(	2857	)	,
(	2858	)	,
(	2859	)	,
(	2860	)	,
(	2861	)	,
(	2862	)	,
(	2863	)	,
(	2864	)	,
(	2864	)	,
(	2865	)	,
(	2866	)	,
(	2867	)	,
(	2868	)	,
(	2869	)	,
(	2870	)	,
(	2871	)	,
(	2872	)	,
(	2873	)	,
(	2874	)	,
(	2874	)	,
(	2875	)	,
(	2876	)	,
(	2877	)	,
(	2878	)	,
(	2879	)	,
(	2880	)	,
(	2881	)	,
(	2882	)	,
(	2883	)	,
(	2884	)	,
(	2885	)	,
(	2886	)	,
(	2886	)	,
(	2887	)	,
(	2888	)	,
(	2889	)	,
(	2890	)	,
(	2891	)	,
(	2892	)	,
(	2893	)	,
(	2894	)	,
(	2895	)	,
(	2896	)	,
(	2897	)	,
(	2898	)	,
(	2899	)	,
(	2899	)	,
(	2900	)	,
(	2901	)	,
(	2902	)	,
(	2903	)	,
(	2904	)	,
(	2905	)	,
(	2906	)	,
(	2907	)	,
(	2908	)	,
(	2909	)	,
(	2910	)	,
(	2911	)	,
(	2912	)	,
(	2913	)	,
(	2914	)	,
(	2915	)	,
(	2915	)	,
(	2916	)	,
(	2917	)	,
(	2918	)	,
(	2919	)	,
(	2920	)	,
(	2921	)	,
(	2922	)	,
(	2923	)	,
(	2924	)	,
(	2925	)	,
(	2926	)	,
(	2927	)	,
(	2928	)	,
(	2929	)	,
(	2930	)	,
(	2931	)	,
(	2932	)	,
(	2933	)	,
(	2934	)	,
(	2934	)	,
(	2935	)	,
(	2936	)	,
(	2937	)	,
(	2938	)	,
(	2939	)	,
(	2940	)	,
(	2941	)	,
(	2942	)	,
(	2943	)	,
(	2944	)	,
(	2945	)	,
(	2946	)	,
(	2947	)	,
(	2948	)	,
(	2949	)	,
(	2950	)	,
(	2951	)	,
(	2952	)	,
(	2953	)	,
(	2954	)	,
(	2955	)	,
(	2956	)	,
(	2957	)	,
(	2958	)	,
(	2959	)	,
(	2960	)	,
(	2961	)	,
(	2962	)	,
(	2962	)	,
(	2963	)	,
(	2964	)	,
(	2965	)	,
(	2966	)	,
(	2967	)	,
(	2968	)	,
(	2969	)	,
(	2970	)	,
(	2971	)	,
(	2972	)	,
(	2973	)	,
(	2974	)	,
(	2975	)	,
(	2976	)	,
(	2977	)	,
(	2978	)	,
(	2979	)	,
(	2980	)	,
(	2981	)	,
(	2982	)	,
(	2983	)	,
(	2984	)	,
(	2985	)	,
(	2986	)	,
(	2987	)	,
(	2988	)	,
(	2989	)	,
(	2990	)	,
(	2991	)	,
(	2992	)	,
(	2993	)	,
(	2994	)	,
(	2995	)	,
(	2996	)	,
(	2997	)	,
(	2998	)	,
(	2999	)	,
(	3000	)	,
(	3001	)	,
(	3002	)	,
(	3003	)	,
(	3004	)	,
(	3005	)	,
(	3006	)	,
(	3007	)	,
(	3008	)	,
(	3009	)	,
(	3010	)	,
(	3011	)	,
(	3012	)	,
(	3013	)	,
(	3014	)	,
(	3015	)	,
(	3016	)	,
(	3017	)	,
(	3018	)	,
(	3019	)	,
(	3020	)	,
(	3021	)	,
(	3022	)	,
(	3023	)	,
(	3024	)	,
(	3025	)	,
(	3026	)	,
(	3027	)	,
(	3028	)	,
(	3029	)	,
(	3030	)	,
(	3031	)	,
(	3032	)	,
(	3033	)	,
(	3034	)	,
(	3035	)	,
(	3036	)	,
(	3037	)	,
(	3038	)	,
(	3040	)	,
(	3041	)	,
(	3042	)	,
(	3043	)	,
(	3044	)	,
(	3045	)	,
(	3046	)	,
(	3047	)	,
(	3048	)	,
(	3049	)	,
(	3050	)	,
(	3051	)	,
(	3052	)	,
(	3053	)	,
(	3054	)	,
(	3055	)	,
(	3056	)	,
(	3057	)	,
(	3058	)	,
(	3059	)	,
(	3060	)	,
(	3061	)	,
(	3062	)	,
(	3063	)	,
(	3064	)	,
(	3065	)	,
(	3066	)	,
(	3067	)	,
(	3069	)	,
(	3070	)	,
(	3071	)	,
(	3072	)	,
(	3073	)	,
(	3074	)	,
(	3075	)	,
(	3076	)	,
(	3077	)	,
(	3078	)	,
(	3079	)	,
(	3080	)	,
(	3081	)	,
(	3082	)	,
(	3083	)	,
(	3084	)	,
(	3085	)	,
(	3086	)	,
(	3087	)	,
(	3089	)	,
(	3090	)	,
(	3091	)	,
(	3092	)	,
(	3093	)	,
(	3094	)	,
(	3095	)	,
(	3096	)	,
(	3097	)	,
(	3098	)	,
(	3099	)	,
(	3100	)	,
(	3101	)	,
(	3102	)	,
(	3103	)	,
(	3105	)	,
(	3106	)	,
(	3107	)	,
(	3108	)	,
(	3109	)	,
(	3110	)	,
(	3111	)	,
(	3112	)	,
(	3113	)	,
(	3114	)	,
(	3115	)	,
(	3116	)	,
(	3117	)	,
(	3119	)	,
(	3120	)	,
(	3121	)	,
(	3122	)	,
(	3123	)	,
(	3124	)	,
(	3125	)	,
(	3126	)	,
(	3127	)	,
(	3128	)	,
(	3129	)	,
(	3130	)	,
(	3132	)	,
(	3133	)	,
(	3134	)	,
(	3135	)	,
(	3136	)	,
(	3137	)	,
(	3138	)	,
(	3139	)	,
(	3140	)	,
(	3141	)	,
(	3142	)	,
(	3144	)	,
(	3145	)	,
(	3146	)	,
(	3147	)	,
(	3148	)	,
(	3149	)	,
(	3150	)	,
(	3151	)	,
(	3152	)	,
(	3153	)	,
(	3155	)	,
(	3156	)	,
(	3157	)	,
(	3158	)	,
(	3159	)	,
(	3160	)	,
(	3161	)	,
(	3162	)	,
(	3163	)	,
(	3165	)	,
(	3166	)	,
(	3167	)	,
(	3168	)	,
(	3169	)	,
(	3170	)	,
(	3171	)	,
(	3172	)	,
(	3173	)	,
(	3175	)	,
(	3176	)	,
(	3177	)	,
(	3178	)	,
(	3179	)	,
(	3180	)	,
(	3181	)	,
(	3182	)	,
(	3184	)	,
(	3185	)	,
(	3186	)	,
(	3187	)	,
(	3188	)	,
(	3189	)	,
(	3190	)	,
(	3191	)	,
(	3193	)	,
(	3194	)	,
(	3195	)	,
(	3196	)	,
(	3197	)	,
(	3198	)	,
(	3199	)	,
(	3201	)	,
(	3202	)	,
(	3203	)	,
(	3204	)	,
(	3205	)	,
(	3206	)	,
(	3207	)	,
(	3209	)	,
(	3210	)	,
(	3211	)	,
(	3212	)	,
(	3213	)	,
(	3214	)	,
(	3215	)	,
(	3217	)	,
(	3218	)	,
(	3219	)	,
(	3220	)	,
(	3221	)	,
(	3222	)	,
(	3223	)	,
(	3225	)	,
(	3226	)	,
(	3227	)	,
(	3228	)	,
(	3229	)	,
(	3230	)	,
(	3232	)	,
(	3233	)	,
(	3234	)	,
(	3235	)	,
(	3236	)	,
(	3237	)	,
(	3239	)	,
(	3240	)	,
(	3241	)	,
(	3242	)	,
(	3243	)	,
(	3244	)	,
(	3246	)	,
(	3247	)	,
(	3248	)	,
(	3249	)	,
(	3250	)	,
(	3251	)	,
(	3253	)	,
(	3254	)	,
(	3255	)	,
(	3256	)	,
(	3257	)	,
(	3259	)	,
(	3260	)	,
(	3261	)	,
(	3262	)	,
(	3263	)	,
(	3264	)	,
(	3266	)	,
(	3267	)	,
(	3268	)	,
(	3269	)	,
(	3270	)	,
(	3272	)	,
(	3273	)	,
(	3274	)	,
(	3275	)	,
(	3276	)	,
(	3277	)	,
(	3279	)	,
(	3280	)	,
(	3281	)	,
(	3282	)	,
(	3283	)	,
(	3285	)	,
(	3286	)	,
(	3287	)	,
(	3288	)	,
(	3289	)	,
(	3291	)	,
(	3292	)	,
(	3293	)	,
(	3294	)	,
(	3295	)	,
(	3297	)	,
(	3298	)	,
(	3299	)	,
(	3300	)	,
(	3302	)	,
(	3303	)	,
(	3304	)	,
(	3305	)	,
(	3306	)	,
(	3308	)	,
(	3309	)	,
(	3310	)	,
(	3311	)	,
(	3312	)	,
(	3314	)	,
(	3315	)	,
(	3316	)	,
(	3317	)	,
(	3319	)	,
(	3320	)	,
(	3321	)	,
(	3322	)	,
(	3323	)	,
(	3325	)	,
(	3326	)	,
(	3327	)	,
(	3328	)	,
(	3330	)	,
(	3331	)	,
(	3332	)	,
(	3333	)	,
(	3335	)	,
(	3336	)	,
(	3337	)	,
(	3338	)	,
(	3340	)	,
(	3341	)	,
(	3342	)	,
(	3343	)	,
(	3344	)	,
(	3346	)	,
(	3347	)	,
(	3348	)	,
(	3349	)	,
(	3351	)	,
(	3352	)	,
(	3353	)	,
(	3354	)	,
(	3356	)	,
(	3357	)	,
(	3358	)	,
(	3359	)	,
(	3361	)	,
(	3362	)	,
(	3363	)	,
(	3364	)	,
(	3366	)	,
(	3367	)	,
(	3368	)	,
(	3370	)	,
(	3371	)	,
(	3372	)	,
(	3373	)	,
(	3375	)	,
(	3376	)	,
(	3377	)	,
(	3378	)	,
(	3380	)	,
(	3381	)	,
(	3382	)	,
(	3383	)	,
(	3385	)	,
(	3386	)	,
(	3387	)	,
(	3389	)	,
(	3390	)	,
(	3391	)	,
(	3392	)	,
(	3394	)	,
(	3395	)	,
(	3396	)	,
(	3398	)	,
(	3399	)	,
(	3400	)	,
(	3401	)	,
(	3403	)	,
(	3404	)	,
(	3405	)	,
(	3407	)	,
(	3408	)	,
(	3409	)	,
(	3410	)	,
(	3412	)	,
(	3413	)	,
(	3414	)	,
(	3416	)	,
(	3417	)	,
(	3418	)	,
(	3419	)	,
(	3421	)	,
(	3422	)	,
(	3423	)	,
(	3425	)	,
(	3426	)	,
(	3427	)	,
(	3429	)	,
(	3430	)	,
(	3431	)	,
(	3432	)	,
(	3434	)	,
(	3435	)	,
(	3436	)	,
(	3438	)	,
(	3439	)	,
(	3440	)	,
(	3442	)	,
(	3443	)	,
(	3444	)	,
(	3446	)	,
(	3447	)	,
(	3448	)	,
(	3450	)	,
(	3451	)	,
(	3452	)	,
(	3454	)	,
(	3455	)	,
(	3456	)	,
(	3458	)	,
(	3459	)	,
(	3460	)	,
(	3462	)	,
(	3463	)	,
(	3464	)	,
(	3466	)	,
(	3467	)	,
(	3468	)	,
(	3470	)	,
(	3471	)	,
(	3472	)	,
(	3474	)	,
(	3475	)	,
(	3476	)	,
(	3478	)	,
(	3479	)	,
(	3480	)	,
(	3482	)	,
(	3483	)	,
(	3484	)	,
(	3486	)	,
(	3487	)	,
(	3488	)	,
(	3490	)	,
(	3491	)	,
(	3492	)	,
(	3494	)	,
(	3495	)	,
(	3497	)	,
(	3498	)	,
(	3499	)	,
(	3501	)	,
(	3502	)	,
(	3503	)	,
(	3505	)	,
(	3506	)	,
(	3507	)	,
(	3509	)	,
(	3510	)	,
(	3512	)	,
(	3513	)	,
(	3514	)	,
(	3516	)	,
(	3517	)	,
(	3518	)	,
(	3520	)	,
(	3521	)	,
(	3523	)	,
(	3524	)	,
(	3525	)	,
(	3527	)	,
(	3528	)	,
(	3529	)	,
(	3531	)	,
(	3532	)	,
(	3534	)	,
(	3535	)	,
(	3536	)	,
(	3538	)	,
(	3539	)	,
(	3541	)	,
(	3542	)	,
(	3543	)	,
(	3545	)	,
(	3546	)	,
(	3547	)	,
(	3549	)	,
(	3550	)	,
(	3552	)	,
(	3553	)	,
(	3555	)	,
(	3556	)	,
(	3557	)	,
(	3559	)	,
(	3560	)	,
(	3562	)	,
(	3563	)	,
(	3564	)	,
(	3566	)	,
(	3567	)	,
(	3569	)	,
(	3570	)	,
(	3571	)	,
(	3573	)	,
(	3574	)	,
(	3576	)	,
(	3577	)	,
(	3579	)	,
(	3580	)	,
(	3581	)	,
(	3583	)	,
(	3584	)	,
(	3586	)	,
(	3587	)	,
(	3589	)	,
(	3590	)	,
(	3591	)	,
(	3593	)	,
(	3594	)	,
(	3596	)	,
(	3597	)	,
(	3599	)	,
(	3600	)	,
(	3601	)	,
(	3603	)	,
(	3604	)	,
(	3606	)	,
(	3607	)	,
(	3609	)	,
(	3610	)	,
(	3612	)	,
(	3613	)	,
(	3614	)	,
(	3616	)	,
(	3617	)	,
(	3619	)	,
(	3620	)	,
(	3622	)	,
(	3623	)	,
(	3625	)	,
(	3626	)	,
(	3628	)	,
(	3629	)	,
(	3630	)	,
(	3632	)	,
(	3633	)	,
(	3635	)	,
(	3636	)	,
(	3638	)	,
(	3639	)	,
(	3641	)	,
(	3642	)	,
(	3644	)	,
(	3645	)	,
(	3647	)	,
(	3648	)	,
(	3650	)	,
(	3651	)	,
(	3653	)	,
(	3654	)	,
(	3656	)	,
(	3657	)	,
(	3659	)	,
(	3660	)	,
(	3662	)	,
(	3663	)	,
(	3664	)	,
(	3666	)	,
(	3667	)	,
(	3669	)	,
(	3670	)	,
(	3672	)	,
(	3673	)	,
(	3675	)	,
(	3676	)	,
(	3678	)	,
(	3679	)	,
(	3681	)	,
(	3682	)	,
(	3684	)	,
(	3686	)	,
(	3687	)	,
(	3689	)	,
(	3690	)	,
(	3692	)	,
(	3693	)	,
(	3695	)	,
(	3696	)	,
(	3698	)	,
(	3699	)	,
(	3701	)	,
(	3702	)	,
(	3704	)	,
(	3705	)	,
(	3707	)	,
(	3708	)	,
(	3710	)	,
(	3711	)	,
(	3713	)	,
(	3714	)	,
(	3716	)	,
(	3717	)	,
(	3719	)	,
(	3721	)	,
(	3722	)	,
(	3724	)	,
(	3725	)	,
(	3727	)	,
(	3728	)	,
(	3730	)	,
(	3731	)	,
(	3733	)	,
(	3734	)	,
(	3736	)	,
(	3738	)	,
(	3739	)	,
(	3741	)	,
(	3742	)	,
(	3744	)	,
(	3745	)	,
(	3747	)	,
(	3748	)	,
(	3750	)	,
(	3752	)	,
(	3753	)	,
(	3755	)	,
(	3756	)	,
(	3758	)	,
(	3759	)	,
(	3761	)	,
(	3763	)	,
(	3764	)	,
(	3766	)	,
(	3767	)	,
(	3769	)	,
(	3770	)	,
(	3772	)	,
(	3774	)	,
(	3775	)	,
(	3777	)	,
(	3778	)	,
(	3780	)	,
(	3782	)	,
(	3783	)	,
(	3785	)	,
(	3786	)	,
(	3788	)	,
(	3789	)	,
(	3791	)	,
(	3793	)	,
(	3794	)	,
(	3796	)	,
(	3797	)	,
(	3799	)	,
(	3801	)	,
(	3802	)	,
(	3804	)	,
(	3805	)	,
(	3807	)	,
(	3809	)	,
(	3810	)	,
(	3812	)	,
(	3814	)	,
(	3815	)	,
(	3817	)	,
(	3818	)	,
(	3820	)	,
(	3822	)	,
(	3823	)	,
(	3825	)	,
(	3827	)	,
(	3828	)	,
(	3830	)	,
(	3831	)	,
(	3833	)	,
(	3835	)	,
(	3836	)	,
(	3838	)	,
(	3840	)	,
(	3841	)	,
(	3843	)	,
(	3845	)	,
(	3846	)	,
(	3848	)	,
(	3849	)	,
(	3851	)	,
(	3853	)	,
(	3854	)	,
(	3856	)	,
(	3858	)	,
(	3859	)	,
(	3861	)	,
(	3863	)	,
(	3864	)	,
(	3866	)	,
(	3868	)	,
(	3869	)	,
(	3871	)	,
(	3873	)	,
(	3874	)	,
(	3876	)	,
(	3878	)	,
(	3879	)	,
(	3881	)	,
(	3883	)	,
(	3884	)	,
(	3886	)	,
(	3888	)	,
(	3889	)	,
(	3891	)	,
(	3893	)	,
(	3894	)	,
(	3896	)	,
(	3898	)	,
(	3899	)	,
(	3901	)	,
(	3903	)	,
(	3905	)	,
(	3906	)	,
(	3908	)	,
(	3910	)	,
(	3911	)	,
(	3913	)	,
(	3915	)	,
(	3916	)	,
(	3918	)	,
(	3920	)	,
(	3922	)	,
(	3923	)	,
(	3925	)	,
(	3927	)	,
(	3928	)	,
(	3930	)	,
(	3932	)	,
(	3934	)	,
(	3935	)	,
(	3937	)	,
(	3939	)	,
(	3940	)	,
(	3942	)	,
(	3944	)	,
(	3946	)	,
(	3947	)	,
(	3949	)	,
(	3951	)	,
(	3953	)	,
(	3954	)	,
(	3956	)	,
(	3958	)	,
(	3960	)	,
(	3961	)	,
(	3963	)	,
(	3965	)	,
(	3967	)	,
(	3968	)	,
(	3970	)	,
(	3972	)	,
(	3974	)	,
(	3975	)	,
(	3977	)	,
(	3979	)	,
(	3981	)	,
(	3982	)	,
(	3984	)	,
(	3986	)	,
(	3988	)	,
(	3989	)	,
(	3991	)	,
(	3993	)	,
(	3995	)	,
(	3996	)	,
(	3998	)	,
(	4000	)	,
(	4002	)	,
(	4004	)	,
(	4005	)	,
(	4007	)	,
(	4009	)	,
(	4011	)	,
(	4012	)	,
(	4014	)	,
(	4016	)	,
(	4018	)	,
(	4020	)	,
(	4021	)	,
(	4023	)	,
(	4025	)	,
(	4027	)	,
(	4029	)	,
(	4030	)	,
(	4032	)	,
(	4034	)	,
(	4036	)	,
(	4038	)	,
(	4039	)	,
(	4041	)	,
(	4043	)	,
(	4045	)	,
(	4047	)	,
(	4049	)	,
(	4050	)	,
(	4052	)	,
(	4054	)	,
(	4056	)	,
(	4058	)	,
(	4060	)	,
(	4061	)	,
(	4063	)	,
(	4065	)	,
(	4067	)	,
(	4069	)	,
(	4071	)	,
(	4072	)	,
(	4074	)	,
(	4076	)	,
(	4078	)	,
(	4080	)	,
(	4082	)	,
(	4083	)	,
(	4085	)	,
(	4087	)	,
(	4089	)	,
(	4091	)	,
(	4093	)	,
(	4095	)	,
(	4096	)	,
(	4098	)	,
(	4100	)	,
(	4102	)	,
(	4104	)	,
(	4106	)	,
(	4108	)	,
(	4110	)	,
(	4111	)	,
(	4113	)	,
(	4115	)	,
(	4117	)	,
(	4119	)	,
(	4121	)	,
(	4123	)	,
(	4125	)	,
(	4127	)	,
(	4128	)	,
(	4130	)	,
(	4132	)	,
(	4134	)	,
(	4136	)	,
(	4138	)	,
(	4140	)	,
(	4142	)	,
(	4144	)	,
(	4146	)	,
(	4147	)	,
(	4149	)	,
(	4151	)	,
(	4153	)	,
(	4155	)	,
(	4157	)	,
(	4159	)	,
(	4161	)	,
(	4163	)	,
(	4165	)	,
(	4167	)	,
(	4169	)	,
(	4171	)	,
(	4172	)	,
(	4174	)	,
(	4176	)	,
(	4178	)	,
(	4180	)	,
(	4182	)	,
(	4184	)	,
(	4186	)	,
(	4188	)	,
(	4190	)	,
(	4192	)	,
(	4194	)	,
(	4196	)	,
(	4198	)	,
(	4200	)	,
(	4202	)	,
(	4204	)	,
(	4206	)	,
(	4208	)	,
(	4210	)	,
(	4212	)	,
(	4213	)	,
(	4215	)	,
(	4217	)	,
(	4219	)	,
(	4221	)	,
(	4223	)	,
(	4225	)	,
(	4227	)	,
(	4229	)	,
(	4231	)	,
(	4233	)	,
(	4235	)	,
(	4237	)	,
(	4239	)	,
(	4241	)	,
(	4243	)	,
(	4245	)	,
(	4247	)	,
(	4249	)	,
(	4251	)	,
(	4253	)	,
(	4255	)	,
(	4257	)	,
(	4259	)	,
(	4261	)	,
(	4263	)	,
(	4265	)	,
(	4267	)	,
(	4269	)	,
(	4271	)	,
(	4274	)	,
(	4276	)	,
(	4278	)	,
(	4280	)	,
(	4282	)	,
(	4284	)	,
(	4286	)	,
(	4288	)	,
(	4290	)	,
(	4292	)	,
(	4294	)	,
(	4296	)	,
(	4298	)	,
(	4300	)	,
(	4302	)	,
(	4304	)	,
(	4306	)	,
(	4308	)	,
(	4310	)	,
(	4312	)	,
(	4314	)	,
(	4317	)	,
(	4319	)	,
(	4321	)	,
(	4323	)	,
(	4325	)	,
(	4327	)	,
(	4329	)	,
(	4331	)	,
(	4333	)	,
(	4335	)	,
(	4337	)	,
(	4339	)	,
(	4342	)	,
(	4344	)	,
(	4346	)	,
(	4348	)	,
(	4350	)	,
(	4352	)	,
(	4354	)	,
(	4356	)	,
(	4358	)	,
(	4360	)	,
(	4363	)	,
(	4365	)	,
(	4367	)	,
(	4369	)	,
(	4371	)	,
(	4373	)	,
(	4375	)	,
(	4377	)	,
(	4380	)	,
(	4382	)	,
(	4384	)	,
(	4386	)	,
(	4388	)	,
(	4390	)	,
(	4392	)	,
(	4395	)	,
(	4397	)	,
(	4399	)	,
(	4401	)	,
(	4403	)	,
(	4405	)	,
(	4407	)	,
(	4410	)	,
(	4412	)	,
(	4414	)	,
(	4416	)	,
(	4418	)	,
(	4420	)	,
(	4423	)	,
(	4425	)	,
(	4427	)	,
(	4429	)	,
(	4431	)	,
(	4433	)	,
(	4436	)	,
(	4438	)	,
(	4440	)	,
(	4442	)	,
(	4444	)	,
(	4447	)	,
(	4449	)	,
(	4451	)	,
(	4453	)	,
(	4455	)	,
(	4458	)	,
(	4460	)	,
(	4462	)	,
(	4464	)	,
(	4467	)	,
(	4469	)	,
(	4471	)	,
(	4473	)	,
(	4475	)	,
(	4478	)	,
(	4480	)	,
(	4482	)	,
(	4484	)	,
(	4487	)	,
(	4489	)	,
(	4491	)	,
(	4493	)	,
(	4496	)	,
(	4498	)	,
(	4500	)	,
(	4502	)	,
(	4505	)	,
(	4507	)	,
(	4509	)	,
(	4511	)	,
(	4514	)	,
(	4516	)	,
(	4518	)	,
(	4520	)	,
(	4523	)	,
(	4525	)	,
(	4527	)	,
(	4529	)	,
(	4532	)	,
(	4534	)	,
(	4536	)	,
(	4539	)	,
(	4541	)	,
(	4543	)	,
(	4545	)	,
(	4548	)	,
(	4550	)	,
(	4552	)	,
(	4555	)	,
(	4557	)	,
(	4559	)	,
(	4562	)	,
(	4564	)	,
(	4566	)	,
(	4569	)	,
(	4571	)	,
(	4573	)	,
(	4575	)	,
(	4578	)	,
(	4580	)	,
(	4582	)	,
(	4585	)	,
(	4587	)	,
(	4589	)	,
(	4592	)	,
(	4594	)	,
(	4597	)	,
(	4599	)	,
(	4601	)	,
(	4604	)	,
(	4606	)	,
(	4608	)	,
(	4611	)	,
(	4613	)	,
(	4615	)	,
(	4618	)	,
(	4620	)	,
(	4622	)	,
(	4625	)	,
(	4627	)	,
(	4630	)	,
(	4632	)	,
(	4634	)	,
(	4637	)	,
(	4639	)	,
(	4642	)	,
(	4644	)	,
(	4646	)	,
(	4649	)	,
(	4651	)	,
(	4654	)	,
(	4656	)	,
(	4658	)	,
(	4661	)	,
(	4663	)	,
(	4666	)	,
(	4668	)	,
(	4670	)	,
(	4673	)	,
(	4675	)	,
(	4678	)	,
(	4680	)	,
(	4683	)	,
(	4685	)	,
(	4688	)	,
(	4690	)	,
(	4692	)	,
(	4695	)	,
(	4697	)	,
(	4700	)	,
(	4702	)	,
(	4705	)	,
(	4707	)	,
(	4710	)	,
(	4712	)	,
(	4715	)	,
(	4717	)	,
(	4719	)	,
(	4722	)	,
(	4724	)	,
(	4727	)	,
(	4729	)	,
(	4732	)	,
(	4734	)	,
(	4737	)	,
(	4739	)	,
(	4742	)	,
(	4744	)	,
(	4747	)	,
(	4749	)	,
(	4752	)	,
(	4754	)	,
(	4757	)	,
(	4759	)	,
(	4762	)	,
(	4764	)	,
(	4767	)	,
(	4769	)	,
(	4772	)	,
(	4775	)	,
(	4777	)	,
(	4780	)	,
(	4782	)	,
(	4785	)	,
(	4787	)	,
(	4790	)	,
(	4792	)	,
(	4795	)	,
(	4797	)	,
(	4800	)	,
(	4803	)	,
(	4805	)	,
(	4808	)	,
(	4810	)	,
(	4813	)	,
(	4815	)	,
(	4818	)	,
(	4821	)	,
(	4823	)	,
(	4826	)	,
(	4828	)	,
(	4831	)	,
(	4834	)	,
(	4836	)	,
(	4839	)	,
(	4841	)	,
(	4844	)	,
(	4847	)	,
(	4849	)	,
(	4852	)	,
(	4854	)	,
(	4857	)	,
(	4860	)	,
(	4862	)	,
(	4865	)	,
(	4867	)	,
(	4870	)	,
(	4873	)	,
(	4875	)	,
(	4878	)	,
(	4881	)	,
(	4883	)	,
(	4886	)	,
(	4889	)	,
(	4891	)	,
(	4894	)	,
(	4897	)	,
(	4899	)	,
(	4902	)	,
(	4905	)	,
(	4907	)	,
(	4910	)	,
(	4913	)	,
(	4915	)	,
(	4918	)	,
(	4921	)	,
(	4923	)	,
(	4926	)	,
(	4929	)	,
(	4932	)	,
(	4934	)	,
(	4937	)	,
(	4940	)	,
(	4942	)	,
(	4945	)	,
(	4948	)	,
(	4950	)	,
(	4953	)	,
(	4956	)	,
(	4959	)	,
(	4961	)	,
(	4964	)	,
(	4967	)	,
(	4970	)	,
(	4972	)	,
(	4975	)	,
(	4978	)	,
(	4981	)	,
(	4983	)	,
(	4986	)	,
(	4989	)	,
(	4992	)	,
(	4994	)	,
(	4997	)	,
(	5000	)	,
(	5003	)	,
(	5006	)	,
(	5008	)	,
(	5011	)	,
(	5014	)	,
(	5017	)	,
(	5020	)	,
(	5022	)	,
(	5025	)	,
(	5028	)	,
(	5031	)	,
(	5034	)	,
(	5036	)	,
(	5039	)	,
(	5042	)	,
(	5045	)	,
(	5048	)	,
(	5051	)	,
(	5053	)	,
(	5056	)	,
(	5059	)	,
(	5062	)	,
(	5065	)	,
(	5068	)	,
(	5070	)	,
(	5073	)	,
(	5076	)	,
(	5079	)	,
(	5082	)	,
(	5085	)	,
(	5088	)	,
(	5090	)	,
(	5093	)	,
(	5096	)	,
(	5099	)	,
(	5102	)	,
(	5105	)	,
(	5108	)	,
(	5111	)	,
(	5114	)	,
(	5117	)	,
(	5119	)	,
(	5122	)	,
(	5125	)	,
(	5128	)	,
(	5131	)	,
(	5134	)	,
(	5137	)	,
(	5140	)	,
(	5143	)	,
(	5146	)	,
(	5149	)	,
(	5152	)	,
(	5155	)	,
(	5158	)	,
(	5161	)	,
(	5164	)	,
(	5166	)	,
(	5169	)	,
(	5172	)	,
(	5175	)	,
(	5178	)	,
(	5181	)	,
(	5184	)	,
(	5187	)	,
(	5190	)	,
(	5193	)	,
(	5196	)	,
(	5199	)	,
(	5202	)	,
(	5205	)	,
(	5208	)	,
(	5211	)	,
(	5214	)	,
(	5217	)	,
(	5220	)	,
(	5223	)	,
(	5226	)	,
(	5230	)	,
(	5233	)	,
(	5236	)	,
(	5239	)	,
(	5242	)	,
(	5245	)	,
(	5248	)	,
(	5251	)	,
(	5254	)	,
(	5257	)	,
(	5260	)	,
(	5263	)	,
(	5266	)	,
(	5269	)	,
(	5272	)	,
(	5275	)	,
(	5279	)	,
(	5282	)	,
(	5285	)	,
(	5288	)	,
(	5291	)	,
(	5294	)	,
(	5297	)	,
(	5300	)	,
(	5303	)	,
(	5307	)	,
(	5310	)	,
(	5313	)	,
(	5316	)	,
(	5319	)	,
(	5322	)	,
(	5325	)	,
(	5329	)	,
(	5332	)	,
(	5335	)	,
(	5338	)	,
(	5341	)	,
(	5344	)	,
(	5348	)	,
(	5351	)	,
(	5354	)	,
(	5357	)	,
(	5360	)	,
(	5364	)	,
(	5367	)	,
(	5370	)	,
(	5373	)	,
(	5376	)	,
(	5380	)	,
(	5383	)	,
(	5386	)	,
(	5389	)	,
(	5392	)	,
(	5396	)	,
(	5399	)	,
(	5402	)	,
(	5405	)	,
(	5409	)	,
(	5412	)	,
(	5415	)	,
(	5418	)	,
(	5422	)	,
(	5425	)	,
(	5428	)	,
(	5432	)	,
(	5435	)	,
(	5438	)	,
(	5441	)	,
(	5445	)	,
(	5448	)	,
(	5451	)	,
(	5455	)	,
(	5458	)	,
(	5461	)	,
(	5464	)	,
(	5468	)	,
(	5471	)	,
(	5474	)	,
(	5478	)	,
(	5481	)	,
(	5484	)	,
(	5488	)	,
(	5491	)	,
(	5495	)	,
(	5498	)	,
(	5501	)	,
(	5505	)	,
(	5508	)	,
(	5511	)	,
(	5515	)	,
(	5518	)	,
(	5521	)	,
(	5525	)	,
(	5528	)	,
(	5532	)	,
(	5535	)	,
(	5538	)	,
(	5542	)	,
(	5545	)	,
(	5549	)	,
(	5552	)	,
(	5556	)	,
(	5559	)	,
(	5562	)	,
(	5566	)	,
(	5569	)	,
(	5573	)	,
(	5576	)	,
(	5580	)	,
(	5583	)	,
(	5587	)	,
(	5590	)	,
(	5594	)	,
(	5597	)	,
(	5600	)	,
(	5604	)	,
(	5607	)	,
(	5611	)	,
(	5614	)	,
(	5618	)	,
(	5621	)	,
(	5625	)	,
(	5629	)	,
(	5632	)	,
(	5636	)	,
(	5639	)	,
(	5643	)	,
(	5646	)	,
(	5650	)	,
(	5653	)	,
(	5657	)	,
(	5660	)	,
(	5664	)	,
(	5668	)	,
(	5671	)	,
(	5675	)	,
(	5678	)	,
(	5682	)	,
(	5685	)	,
(	5689	)	,
(	5693	)	,
(	5696	)	,
(	5700	)	,
(	5703	)	,
(	5707	)	,
(	5711	)	,
(	5714	)	,
(	5718	)	,
(	5722	)	,
(	5725	)	,
(	5729	)	,
(	5732	)	,
(	5736	)	,
(	5740	)	,
(	5743	)	,
(	5747	)	,
(	5751	)	,
(	5754	)	,
(	5758	)	,
(	5762	)	,
(	5766	)	,
(	5769	)	,
(	5773	)	,
(	5777	)	,
(	5780	)	,
(	5784	)	,
(	5788	)	,
(	5792	)	,
(	5795	)	,
(	5799	)	,
(	5803	)	,
(	5806	)	,
(	5810	)	,
(	5814	)	,
(	5818	)	,
(	5821	)	,
(	5825	)	,
(	5829	)	,
(	5833	)	,
(	5837	)	,
(	5840	)	,
(	5844	)	,
(	5848	)	,
(	5852	)	,
(	5856	)	,
(	5859	)	,
(	5863	)	,
(	5867	)	,
(	5871	)	,
(	5875	)	,
(	5879	)	,
(	5882	)	,
(	5886	)	,
(	5890	)	,
(	5894	)	,
(	5898	)	,
(	5902	)	,
(	5906	)	,
(	5909	)	,
(	5913	)	,
(	5917	)	,
(	5921	)	,
(	5925	)	,
(	5929	)	,
(	5933	)	,
(	5937	)	,
(	5941	)	,
(	5945	)	,
(	5948	)	,
(	5952	)	,
(	5956	)	,
(	5960	)	,
(	5964	)	,
(	5968	)	,
(	5972	)	,
(	5976	)	,
(	5980	)	,
(	5984	)	,
(	5988	)	,
(	5992	)	,
(	5996	)	,
(	6000	)	,
(	6004	)	,
(	6008	)	,
(	6012	)	,
(	6016	)	,
(	6020	)	,
(	6024	)	,
(	6028	)	,
(	6032	)	,
(	6036	)	,
(	6040	)	,
(	6044	)	,
(	6048	)	,
(	6052	)	,
(	6057	)	,
(	6061	)	,
(	6065	)	,
(	6069	)	,
(	6073	)	,
(	6077	)	,
(	6081	)	,
(	6085	)	,
(	6089	)	,
(	6093	)	,
(	6098	)	,
(	6102	)	,
(	6106	)	,
(	6110	)	,
(	6114	)	,
(	6118	)	,
(	6122	)	,
(	6127	)	,
(	6131	)	,
(	6135	)	,
(	6139	)	,
(	6143	)	,
(	6148	)	,
(	6152	)	,
(	6156	)	,
(	6160	)	,
(	6164	)	,
(	6169	)	,
(	6173	)	,
(	6177	)	,
(	6181	)	,
(	6186	)	,
(	6190	)	,
(	6194	)	,
(	6198	)	,
(	6203	)	,
(	6207	)	,
(	6211	)	,
(	6215	)	,
(	6220	)	,
(	6224	)	,
(	6228	)	,
(	6233	)	,
(	6237	)	,
(	6241	)	,
(	6246	)	,
(	6250	)	,
(	6254	)	,
(	6259	)	,
(	6263	)	,
(	6267	)	,
(	6272	)	,
(	6276	)	,
(	6281	)	,
(	6285	)	,
(	6289	)	,
(	6294	)	,
(	6298	)	,
(	6303	)	,
(	6307	)	,
(	6311	)	,
(	6316	)	,
(	6320	)	,
(	6325	)	,
(	6329	)	,
(	6334	)	,
(	6338	)	,
(	6342	)	,
(	6347	)	,
(	6351	)	,
(	6356	)	,
(	6360	)	,
(	6365	)	,
(	6369	)	,
(	6374	)	,
(	6378	)	,
(	6383	)	,
(	6388	)	,
(	6392	)	,
(	6397	)	,
(	6401	)	,
(	6406	)	,
(	6410	)	,
(	6415	)	,
(	6419	)	,
(	6424	)	,
(	6429	)	,
(	6433	)	,
(	6438	)	,
(	6442	)	,
(	6447	)	,
(	6452	)	,
(	6456	)	,
(	6461	)	,
(	6466	)	,
(	6470	)	,
(	6475	)	,
(	6479	)	,
(	6484	)	,
(	6489	)	,
(	6494	)	,
(	6498	)	,
(	6503	)	,
(	6508	)	,
(	6512	)	,
(	6517	)	,
(	6522	)	,
(	6526	)	,
(	6531	)	,
(	6536	)	,
(	6541	)	,
(	6545	)	,
(	6550	)	,
(	6555	)	,
(	6560	)	,
(	6565	)	,
(	6569	)	,
(	6574	)	,
(	6579	)	,
(	6584	)	,
(	6589	)	,
(	6593	)	,
(	6598	)	,
(	6603	)	,
(	6608	)	,
(	6613	)	,
(	6618	)	,
(	6623	)	,
(	6627	)	,
(	6632	)	,
(	6637	)	,
(	6642	)	,
(	6647	)	,
(	6652	)	,
(	6657	)	,
(	6662	)	,
(	6667	)	,
(	6672	)	,
(	6677	)	,
(	6682	)	,
(	6686	)	,
(	6691	)	,
(	6696	)	,
(	6701	)	,
(	6706	)	,
(	6711	)	,
(	6716	)	,
(	6721	)	,
(	6726	)	,
(	6731	)	,
(	6737	)	,
(	6742	)	,
(	6747	)	,
(	6752	)	,
(	6757	)	,
(	6762	)	,
(	6767	)	,
(	6772	)	,
(	6777	)	,
(	6782	)	,
(	6787	)	,
(	6792	)	,
(	6798	)	,
(	6803	)	,
(	6808	)	,
(	6813	)	,
(	6818	)	,
(	6823	)	,
(	6829	)	,
(	6834	)	,
(	6839	)	,
(	6844	)	,
(	6849	)	,
(	6855	)	,
(	6860	)	,
(	6865	)	,
(	6870	)	,
(	6875	)	,
(	6881	)	,
(	6886	)	,
(	6891	)	,
(	6897	)	,
(	6902	)	,
(	6907	)	,
(	6912	)	,
(	6918	)	,
(	6923	)	,
(	6928	)	,
(	6934	)	,
(	6939	)	,
(	6944	)	,
(	6950	)	,
(	6955	)	,
(	6961	)	,
(	6966	)	,
(	6971	)	,
(	6977	)	,
(	6982	)	,
(	6988	)	,
(	6993	)	,
(	6998	)	,
(	7004	)	,
(	7009	)	,
(	7015	)	,
(	7020	)	,
(	7026	)	,
(	7031	)	,
(	7037	)	,
(	7042	)	,
(	7048	)	,
(	7053	)	,
(	7059	)	,
(	7064	)	,
(	7070	)	,
(	7075	)	,
(	7081	)	,
(	7087	)	,
(	7092	)	,
(	7098	)	,
(	7103	)	,
(	7109	)	,
(	7115	)	,
(	7120	)	,
(	7126	)	,
(	7132	)	,
(	7137	)	,
(	7143	)	,
(	7149	)	,
(	7154	)	,
(	7160	)	,
(	7166	)	,
(	7171	)	,
(	7177	)	,
(	7183	)	,
(	7188	)	,
(	7194	)	,
(	7200	)	,
(	7206	)	,
(	7212	)	,
(	7217	)	,
(	7223	)	,
(	7229	)	,
(	7235	)	,
(	7241	)	,
(	7246	)	,
(	7252	)	,
(	7258	)	,
(	7264	)	,
(	7270	)	,
(	7276	)	,
(	7282	)	,
(	7287	)	,
(	7293	)	,
(	7299	)	,
(	7305	)	,
(	7311	)	,
(	7317	)	,
(	7323	)	,
(	7329	)	,
(	7335	)	,
(	7341	)	,
(	7347	)	,
(	7353	)	,
(	7359	)	,
(	7365	)	,
(	7371	)	,
(	7377	)	,
(	7383	)	,
(	7389	)	,
(	7395	)	,
(	7401	)	,
(	7407	)	,
(	7414	)	,
(	7420	)	,
(	7426	)	,
(	7432	)	,
(	7438	)	,
(	7444	)	,
(	7450	)	,
(	7457	)	,
(	7463	)	,
(	7469	)	,
(	7475	)	,
(	7481	)	,
(	7488	)	,
(	7494	)	,
(	7500	)	,
(	7506	)	,
(	7513	)	,
(	7519	)	,
(	7525	)	,
(	7531	)	,
(	7538	)	,
(	7544	)	,
(	7550	)	,
(	7557	)	,
(	7563	)	,
(	7569	)	,
(	7576	)	,
(	7582	)	,
(	7589	)	,
(	7595	)	,
(	7601	)	,
(	7608	)	,
(	7614	)	,
(	7621	)	,
(	7627	)	,
(	7634	)	,
(	7640	)	,
(	7647	)	,
(	7653	)	,
(	7660	)	,
(	7666	)	,
(	7673	)	,
(	7679	)	,
(	7686	)	,
(	7692	)	,
(	7699	)	,
(	7705	)	,
(	7712	)	,
(	7719	)	,
(	7725	)	,
(	7732	)	,
(	7739	)	,
(	7745	)	,
(	7752	)	,
(	7759	)	,
(	7765	)	,
(	7772	)	,
(	7779	)	,
(	7785	)	,
(	7792	)	,
(	7799	)	,
(	7806	)	,
(	7813	)	,
(	7819	)	,
(	7826	)	,
(	7833	)	,
(	7840	)	,
(	7847	)	,
(	7853	)	,
(	7860	)	,
(	7867	)	,
(	7874	)	,
(	7881	)	,
(	7888	)	,
(	7895	)	,
(	7902	)	,
(	7909	)	,
(	7916	)	,
(	7923	)	,
(	7930	)	,
(	7937	)	,
(	7944	)	,
(	7951	)	,
(	7958	)	,
(	7965	)	,
(	7972	)	,
(	7979	)	,
(	7986	)	,
(	7993	)	,
(	8000	)	,
(	8007	)	,
(	8014	)	,
(	8021	)	,
(	8029	)	,
(	8036	)	,
(	8043	)	,
(	8050	)	,
(	8057	)	,
(	8065	)	,
(	8072	)	,
(	8079	)	,
(	8086	)	,
(	8094	)	,
(	8101	)	,
(	8108	)	,
(	8115	)	,
(	8123	)	,
(	8130	)	,
(	8137	)	,
(	8145	)	,
(	8152	)	,
(	8160	)	,
(	8167	)	,
(	8174	)	,
(	8182	)	,
(	8189	)	,
(	8197	)	,
(	8204	)	,
(	8212	)	,
(	8219	)	,
(	8227	)	,
(	8234	)	,
(	8242	)	,
(	8249	)	,
(	8257	)	,
(	8264	)	,
(	8272	)	,
(	8280	)	,
(	8287	)	,
(	8295	)	,
(	8303	)	,
(	8310	)	,
(	8318	)	,
(	8326	)	,
(	8333	)	,
(	8341	)	,
(	8349	)	,
(	8357	)	,
(	8364	)	,
(	8372	)	,
(	8380	)	,
(	8388	)	,
(	8396	)	,
(	8403	)	,
(	8411	)	,
(	8419	)	,
(	8427	)	,
(	8435	)	,
(	8443	)	,
(	8451	)	,
(	8459	)	,
(	8467	)	,
(	8475	)	,
(	8483	)	,
(	8491	)	,
(	8499	)	,
(	8507	)	,
(	8515	)	,
(	8523	)	,
(	8531	)	,
(	8539	)	,
(	8547	)	,
(	8555	)	,
(	8563	)	,
(	8571	)	,
(	8580	)	,
(	8588	)	,
(	8596	)	,
(	8604	)	,
(	8612	)	,
(	8621	)	,
(	8629	)	,
(	8637	)	,
(	8646	)	,
(	8654	)	,
(	8662	)	,
(	8671	)	,
(	8679	)	,
(	8687	)	,
(	8696	)	,
(	8704	)	,
(	8712	)	,
(	8721	)	,
(	8729	)	,
(	8738	)	,
(	8746	)	,
(	8755	)	,
(	8763	)	,
(	8772	)	,
(	8780	)	,
(	8789	)	,
(	8798	)	,
(	8806	)	,
(	8815	)	,
(	8824	)	,
(	8832	)	,
(	8841	)	,
(	8850	)	,
(	8858	)	,
(	8867	)	,
(	8876	)	,
(	8885	)	,
(	8893	)	,
(	8902	)	,
(	8911	)	,
(	8920	)	,
(	8929	)	,
(	8937	)	,
(	8946	)	,
(	8955	)	,
(	8964	)	,
(	8973	)	,
(	8982	)	,
(	8991	)	,
(	9000	)	,
(	9009	)	,
(	9018	)	,
(	9027	)	,
(	9036	)	,
(	9045	)	,
(	9054	)	,
(	9063	)	,
(	9073	)	,
(	9082	)	,
(	9091	)	,
(	9100	)	,
(	9109	)	,
(	9119	)	,
(	9128	)	,
(	9137	)	,
(	9146	)	,
(	9156	)	,
(	9165	)	,
(	9174	)	,
(	9184	)	,
(	9193	)	,
(	9202	)	,
(	9212	)	,
(	9221	)	,
(	9231	)	,
(	9240	)	,
(	9250	)	,
(	9259	)	,
(	9269	)	,
(	9278	)	,
(	9288	)	,
(	9298	)	,
(	9307	)	,
(	9317	)	,
(	9326	)	,
(	9336	)	,
(	9346	)	,
(	9356	)	,
(	9365	)	,
(	9375	)	,
(	9385	)	,
(	9395	)	,
(	9404	)	,
(	9414	)	,
(	9424	)	,
(	9434	)	,
(	9444	)	,
(	9454	)	,
(	9464	)	,
(	9474	)	,
(	9484	)	,
(	9494	)	,
(	9504	)	,
(	9514	)	,
(	9524	)	,
(	9534	)	,
(	9544	)	,
(	9554	)	,
(	9564	)	,
(	9574	)	,
(	9585	)	,
(	9595	)	,
(	9605	)	,
(	9615	)	,
(	9626	)	,
(	9636	)	,
(	9646	)	,
(	9657	)	,
(	9667	)	,
(	9677	)	,
(	9688	)	,
(	9698	)	,
(	9709	)	,
(	9719	)	,
(	9730	)	,
(	9740	)	,
(	9751	)	,
(	9761	)	,
(	9772	)	,
(	9783	)	,
(	9793	)	,
(	9804	)	,
(	9815	)	,
(	9825	)	,
(	9836	)	,
(	9847	)	,
(	9858	)	,
(	9868	)	,
(	9879	)	,
(	9890	)	,
(	9901	)	,
(	9912	)	,
(	9923	)	,
(	9934	)	,
(	9945	)	,
(	9956	)	,
(	9967	)	,
(	9978	)	,
(	9989	)	,
(	10000	)	,
(	10011	)	,
(	10022	)	,
(	10033	)	,
(	10045	)	,
(	10056	)	,
(	10067	)	,
(	10078	)	,
(	10090	)	,
(	10101	)	,
(	10112	)	,
(	10124	)	,
(	10135	)	,
(	10147	)	,
(	10158	)	,
(	10169	)	,
(	10181	)	,
(	10193	)	,
(	10204	)	,
(	10216	)	,
(	10227	)	,
(	10239	)	,
(	10251	)	,
(	10262	)	,
(	10274	)	,
(	10286	)	,
(	10297	)	,
(	10309	)	,
(	10321	)	,
(	10333	)	,
(	10345	)	,
(	10357	)	,
(	10369	)	,
(	10381	)	,
(	10393	)	,
(	10405	)	,
(	10417	)	,
(	10429	)	,
(	10441	)	,
(	10453	)	,
(	10465	)	,
(	10477	)	,
(	10490	)	,
(	10502	)	,
(	10514	)	,
(	10526	)	,
(	10539	)	,
(	10551	)	,
(	10563	)	,
(	10576	)	,
(	10588	)	,
(	10601	)	,
(	10613	)	,
(	10626	)	,
(	10638	)	,
(	10651	)	,
(	10664	)	,
(	10676	)	,
(	10689	)	,
(	10702	)	,
(	10714	)	,
(	10727	)	,
(	10740	)	,
(	10753	)	,
(	10766	)	,
(	10778	)	,
(	10791	)	,
(	10804	)	,
(	10817	)	,
(	10830	)	,
(	10843	)	,
(	10856	)	,
(	10870	)	,
(	10883	)	,
(	10896	)	,
(	10909	)	,
(	10922	)	,
(	10936	)	,
(	10949	)	,
(	10962	)	,
(	10976	)	,
(	10989	)	,
(	11002	)	,
(	11016	)	,
(	11029	)	,
(	11043	)	,
(	11057	)	,
(	11070	)	,
(	11084	)	,
(	11097	)	,
(	11111	)	,
(	11125	)	,
(	11139	)	,
(	11152	)	,
(	11166	)	,
(	11180	)	,
(	11194	)	,
(	11208	)	,
(	11222	)	,
(	11236	)	,
(	11250	)	,
(	11264	)	,
(	11278	)	,
(	11292	)	,
(	11307	)	,
(	11321	)	,
(	11335	)	,
(	11349	)	,
(	11364	)	,
(	11378	)	,
(	11392	)	,
(	11407	)	,
(	11421	)	,
(	11436	)	,
(	11450	)	,
(	11465	)	,
(	11480	)	,
(	11494	)	,
(	11509	)	,
(	11524	)	,
(	11538	)	,
(	11553	)	,
(	11568	)	,
(	11583	)	,
(	11598	)	,
(	11613	)	,
(	11628	)	,
(	11643	)	,
(	11658	)	,
(	11673	)	,
(	11688	)	,
(	11704	)	,
(	11719	)	,
(	11734	)	,
(	11749	)	,
(	11765	)	,
(	11780	)	,
(	11796	)	,
(	11811	)	,
(	11827	)	,
(	11842	)	,
(	11858	)	,
(	11873	)	,
(	11889	)	,
(	11905	)	,
(	11921	)	,
(	11936	)	,
(	11952	)	,
(	11968	)	,
(	11984	)	,
(	12000	)	,
(	12016	)	,
(	12032	)	,
(	12048	)	,
(	12064	)	,
(	12081	)	,
(	12097	)	,
(	12113	)	,
(	12129	)	,
(	12146	)	,
(	12162	)	,
(	12179	)	,
(	12195	)	,
(	12212	)	,
(	12228	)	,
(	12245	)	,
(	12262	)	,
(	12278	)	,
(	12295	)	,
(	12312	)	,
(	12329	)	,
(	12346	)	,
(	12363	)	,
(	12380	)	,
(	12397	)	,
(	12414	)	,
(	12431	)	,
(	12448	)	,
(	12465	)	,
(	12483	)	,
(	12500	)	,
(	12517	)	,
(	12535	)	,
(	12552	)	,
(	12570	)	,
(	12587	)	,
(	12605	)	,
(	12623	)	,
(	12640	)	,
(	12658	)	,
(	12676	)	,
(	12694	)	,
(	12712	)	,
(	12730	)	,
(	12748	)	,
(	12766	)	,
(	12784	)	,
(	12802	)	,
(	12821	)	,
(	12839	)	,
(	12857	)	,
(	12876	)	,
(	12894	)	,
(	12912	)	,
(	12931	)	,
(	12950	)	,
(	12968	)	,
(	12987	)	,
(	13006	)	,
(	13025	)	,
(	13043	)	,
(	13062	)	,
(	13081	)	,
(	13100	)	,
(	13120	)	,
(	13139	)	,
(	13158	)	,
(	13177	)	,
(	13196	)	,
(	13216	)	,
(	13235	)	,
(	13255	)	,
(	13274	)	,
(	13294	)	,
(	13314	)	,
(	13333	)	,
(	13353	)	,
(	13373	)	,
(	13393	)	,
(	13413	)	,
(	13433	)	,
(	13453	)	,
(	13473	)	,
(	13493	)	,
(	13514	)	,
(	13534	)	,
(	13554	)	,
(	13575	)	,
(	13595	)	,
(	13616	)	,
(	13636	)	,
(	13657	)	,
(	13678	)	,
(	13699	)	,
(	13720	)	,
(	13740	)	,
(	13761	)	,
(	13783	)	,
(	13804	)	,
(	13825	)	,
(	13846	)	,
(	13867	)	,
(	13889	)	,
(	13910	)	,
(	13932	)	,
(	13953	)	,
(	13975	)	,
(	13997	)	,
(	14019	)	,
(	14041	)	,
(	14063	)	,
(	14085	)	,
(	14107	)	,
(	14129	)	,
(	14151	)	,
(	14173	)	,
(	14196	)	,
(	14218	)	,
(	14241	)	,
(	14263	)	,
(	14286	)	,
(	14308	)	,
(	14331	)	,
(	14354	)	,
(	14377	)	,
(	14400	)	,
(	14423	)	,
(	14446	)	,
(	14469	)	,
(	14493	)	,
(	14516	)	,
(	14540	)	,
(	14563	)	,
(	14587	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	,
(	0	)	







);


begin
   -- This is the only statement required. It looks up the converted value of 
	-- the voltage input (in mV) in the v2d_LUT look-up table, and outputs the 
	-- distance (in 10^-4 m) in std_logic_vector format.
    	
   frequency <= std_logic_vector(to_unsigned(v2d_LUT(to_integer(unsigned(voltage))),frequency'length));
	
end behavior;
